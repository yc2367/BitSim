`ifndef __vert_32_tb_V__
`define __vert_32_tb_V__

`include "mac_unit_Vert_32_no_mul.v"

module vert_32_tb;
    
    parameter DATA_WIDTH    = 8;
    parameter VEC_LENGTH    = 32;
    parameter MUX_SEL_WIDTH = 3;
    parameter SUM_ACT_WIDTH = $clog2(VEC_LENGTH) + DATA_WIDTH - 2;
    parameter ACC_WIDTH     = DATA_WIDTH + 16;
    parameter RESULT_WIDTH  = 2*DATA_WIDTH;

    logic                               clk;
	logic                               reset;
	logic                               en_acc;
	logic                               load_accum;

	logic signed   [DATA_WIDTH-1:0]     act_in   [VEC_LENGTH-1:0];   // input activation (signed)
	logic          [MUX_SEL_WIDTH-1:0]  act_sel_in  [VEC_LENGTH/2-1:0]; // input activation MUX select signal
	logic                               act_val_in  [VEC_LENGTH/2-1:0]; // whether activation is valid
	logic signed   [SUM_ACT_WIDTH-1:0]  sum_act  [VEC_LENGTH/8-1:0]; // sum of a group of activations (signed)

	logic          [2:0]                column_idx;    // current column index for shifting 
	logic                               is_msb;        // specify if the current column is MSB
	logic                               is_skip_zero [VEC_LENGTH/8-1:0];  // specify if skip bit 0
	
	logic signed   [ACC_WIDTH-1:0]      accum_prev;
    logic signed   [RESULT_WIDTH-1:0]   result;

    mac_unit_Vert_32_no_mul_clk #(DATA_WIDTH, VEC_LENGTH, MUX_SEL_WIDTH, SUM_ACT_WIDTH, ACC_WIDTH) s (.*);

  initial
    $monitor ("out=%b", result);

  initial begin
    #0 clk = 0; reset = 1;  en_acc = 0;
    #1.2 reset = 0; en_acc = 1; load_accum = 0; accum_prev = 0;

    #1 is_msb=1; column_idx=7; act[0] = -26; act[1] = 25; act[2] = -60; act[3] = -120; act[4] = 25; act[5] = 75; act[6] = 116; act[7] = -117; act[8] = -113; act[9] = 118; act[10] = -56; act[11] = -79; act[12] = 54; act[13] = -105; act[14] = -92; act[15] = -90; act[16] = -121; act[17] = 6; act[18] = 19; act[19] = 23; act[20] = -24; act[21] = -104; act[22] = 71; act[23] = -85; act[24] = 10; act[25] = -95; act[26] = 84; act[27] = 10; act[28] = -80; act[29] = -38; act[30] = 68; act[31] = -82; 
    act_sel_in[0] = 3; act_sel_in[1] = 1; act_sel_in[2] = 0; act_sel_in[3] = 1; act_sel_in[4] = 3; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 3; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 3; act_sel_in[11] = 4; act_sel_in[12] = 1; act_sel_in[13] = 4; act_sel_in[14] = 3; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 1; act_sel_in[3] = 4; act_sel_in[4] = 1; act_sel_in[5] = 0; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 0; act_sel_in[13] = 2; act_sel_in[14] = 1; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=5; act_sel_in[0] = 2; act_sel_in[1] = 0; act_sel_in[2] = 2; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 1; act_sel_in[6] = 2; act_sel_in[7] = 4; act_sel_in[8] = 4; act_sel_in[9] = 0; act_sel_in[10] = 0; act_sel_in[11] = 3; act_sel_in[12] = 2; act_sel_in[13] = 2; act_sel_in[14] = 0; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=4; act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 3; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 3; act_sel_in[7] = 2; act_sel_in[8] = 0; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 0; act_sel_in[12] = 4; act_sel_in[13] = 3; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=3; act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 4; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 0; act_sel_in[7] = 1; act_sel_in[8] = 4; act_sel_in[9] = 2; act_sel_in[10] = 2; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=2; act_sel_in[0] = 1; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 4; act_sel_in[4] = 2; act_sel_in[5] = 1; act_sel_in[6] = 1; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 4; act_sel_in[11] = 4; act_sel_in[12] = 3; act_sel_in[13] = 1; act_sel_in[14] = 3; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 2; act_sel_in[1] = 2; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 0; act_sel_in[5] = 0; act_sel_in[6] = 0; act_sel_in[7] = 3; act_sel_in[8] = 4; act_sel_in[9] = 0; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 0; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=0; act_sel_in[0] = 0; act_sel_in[1] = 3; act_sel_in[2] = 1; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 2; act_sel_in[10] = 3; act_sel_in[11] = 1; act_sel_in[12] = 2; act_sel_in[13] = 0; act_sel_in[14] = 2; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 


    #1 is_msb=1; column_idx=7; act[0] = 8; act[1] = -20; act[2] = 103; act[3] = -31; act[4] = -16; act[5] = -34; act[6] = 101; act[7] = -18; act[8] = 115; act[9] = -85; act[10] = -1; act[11] = 99; act[12] = 112; act[13] = 120; act[14] = -47; act[15] = -81; act[16] = -126; act[17] = -72; act[18] = 66; act[19] = -66; act[20] = 20; act[21] = -83; act[22] = -72; act[23] = 58; act[24] = -78; act[25] = -102; act[26] = 106; act[27] = -74; act[28] = -75; act[29] = -40; act[30] = 73; act[31] = -65; 
    act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 1; act_sel_in[5] = 4; act_sel_in[6] = 4; act_sel_in[7] = 3; act_sel_in[8] = 3; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 3; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 3; act_sel_in[1] = 0; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 1; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 3; act_sel_in[12] = 0; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=5; act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 0; act_sel_in[3] = 0; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 3; act_sel_in[11] = 3; act_sel_in[12] = 3; act_sel_in[13] = 3; act_sel_in[14] = 1; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=4; act_sel_in[0] = 2; act_sel_in[1] = 0; act_sel_in[2] = 4; act_sel_in[3] = 3; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 3; act_sel_in[7] = 1; act_sel_in[8] = 2; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 3; act_sel_in[12] = 2; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 1; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 1; act_sel_in[6] = 3; act_sel_in[7] = 0; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 2; act_sel_in[11] = 4; act_sel_in[12] = 3; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=2; act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 3; act_sel_in[3] = 4; act_sel_in[4] = 2; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 2; act_sel_in[10] = 1; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 1; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 2; act_sel_in[1] = 4; act_sel_in[2] = 0; act_sel_in[3] = 1; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 2; act_sel_in[10] = 0; act_sel_in[11] = 0; act_sel_in[12] = 4; act_sel_in[13] = 3; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 2; act_sel_in[1] = 2; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 0; act_sel_in[7] = 4; act_sel_in[8] = 2; act_sel_in[9] = 3; act_sel_in[10] = 1; act_sel_in[11] = 3; act_sel_in[12] = 1; act_sel_in[13] = 0; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 


    #1 is_msb=1; column_idx=7; act[0] = -126; act[1] = 119; act[2] = 78; act[3] = -97; act[4] = 123; act[5] = 117; act[6] = -1; act[7] = -48; act[8] = -115; act[9] = -17; act[10] = -90; act[11] = 41; act[12] = -73; act[13] = -85; act[14] = -37; act[15] = -124; act[16] = 115; act[17] = -90; act[18] = -70; act[19] = -122; act[20] = -29; act[21] = 34; act[22] = -36; act[23] = 122; act[24] = 47; act[25] = -43; act[26] = -75; act[27] = -36; act[28] = 94; act[29] = 55; act[30] = 30; act[31] = 48; 
    act_sel_in[0] = 4; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 2; act_sel_in[4] = 3; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 2; act_sel_in[11] = 2; act_sel_in[12] = 0; act_sel_in[13] = 4; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 4; act_sel_in[1] = 3; act_sel_in[2] = 1; act_sel_in[3] = 3; act_sel_in[4] = 0; act_sel_in[5] = 0; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 1; act_sel_in[9] = 2; act_sel_in[10] = 1; act_sel_in[11] = 3; act_sel_in[12] = 1; act_sel_in[13] = 0; act_sel_in[14] = 0; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=5; act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 0; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 1; act_sel_in[9] = 0; act_sel_in[10] = 0; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 3; act_sel_in[14] = 1; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=4; act_sel_in[0] = 4; act_sel_in[1] = 0; act_sel_in[2] = 4; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 4; act_sel_in[1] = 0; act_sel_in[2] = 4; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 4; act_sel_in[6] = 4; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 2; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 0; act_sel_in[14] = 3; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=2; act_sel_in[0] = 0; act_sel_in[1] = 0; act_sel_in[2] = 0; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 4; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 2; act_sel_in[9] = 3; act_sel_in[10] = 1; act_sel_in[11] = 0; act_sel_in[12] = 4; act_sel_in[13] = 1; act_sel_in[14] = 3; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 3; act_sel_in[1] = 1; act_sel_in[2] = 4; act_sel_in[3] = 0; act_sel_in[4] = 2; act_sel_in[5] = 3; act_sel_in[6] = 0; act_sel_in[7] = 2; act_sel_in[8] = 1; act_sel_in[9] = 1; act_sel_in[10] = 4; act_sel_in[11] = 4; act_sel_in[12] = 1; act_sel_in[13] = 4; act_sel_in[14] = 1; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 0; act_sel_in[1] = 0; act_sel_in[2] = 2; act_sel_in[3] = 1; act_sel_in[4] = 0; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 2; act_sel_in[8] = 3; act_sel_in[9] = 4; act_sel_in[10] = 4; act_sel_in[11] = 2; act_sel_in[12] = 0; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 


    #1 is_msb=1; column_idx=7; act[0] = 59; act[1] = 103; act[2] = 12; act[3] = -111; act[4] = 98; act[5] = 29; act[6] = -87; act[7] = 21; act[8] = 25; act[9] = 37; act[10] = -88; act[11] = 45; act[12] = 123; act[13] = 44; act[14] = 63; act[15] = 22; act[16] = -43; act[17] = 118; act[18] = 61; act[19] = -33; act[20] = -124; act[21] = 23; act[22] = 15; act[23] = -118; act[24] = 112; act[25] = 95; act[26] = 95; act[27] = 30; act[28] = -115; act[29] = 4; act[30] = 65; act[31] = -58; 
    act_sel_in[0] = 4; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 2; act_sel_in[4] = 4; act_sel_in[5] = 4; act_sel_in[6] = 3; act_sel_in[7] = 1; act_sel_in[8] = 0; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 3; act_sel_in[12] = 3; act_sel_in[13] = 1; act_sel_in[14] = 1; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 3; act_sel_in[1] = 0; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 4; act_sel_in[9] = 0; act_sel_in[10] = 1; act_sel_in[11] = 1; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=5; act_sel_in[0] = 0; act_sel_in[1] = 0; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 1; act_sel_in[8] = 1; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 3; act_sel_in[12] = 3; act_sel_in[13] = 0; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=4; act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 2; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 1; act_sel_in[10] = 1; act_sel_in[11] = 1; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 1; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 1; act_sel_in[1] = 0; act_sel_in[2] = 2; act_sel_in[3] = 3; act_sel_in[4] = 3; act_sel_in[5] = 0; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 2; act_sel_in[11] = 3; act_sel_in[12] = 3; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=2; act_sel_in[0] = 1; act_sel_in[1] = 0; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 0; act_sel_in[5] = 3; act_sel_in[6] = 0; act_sel_in[7] = 2; act_sel_in[8] = 0; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 3; act_sel_in[12] = 1; act_sel_in[13] = 4; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=1; act_sel_in[0] = 2; act_sel_in[1] = 4; act_sel_in[2] = 0; act_sel_in[3] = 0; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 3; act_sel_in[11] = 2; act_sel_in[12] = 3; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=0; act_sel_in[0] = 1; act_sel_in[1] = 1; act_sel_in[2] = 4; act_sel_in[3] = 1; act_sel_in[4] = 0; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 0; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 3; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 1; act_sel_in[14] = 0; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 


    #1 is_msb=1; column_idx=7; act[0] = 121; act[1] = 106; act[2] = -34; act[3] = -26; act[4] = 79; act[5] = 24; act[6] = 81; act[7] = 76; act[8] = -26; act[9] = 89; act[10] = 92; act[11] = 24; act[12] = -119; act[13] = -92; act[14] = -18; act[15] = 86; act[16] = -125; act[17] = -18; act[18] = -92; act[19] = -42; act[20] = 105; act[21] = -84; act[22] = -21; act[23] = 13; act[24] = -108; act[25] = 120; act[26] = -85; act[27] = 111; act[28] = 93; act[29] = 126; act[30] = 105; act[31] = 59; 
    act_sel_in[0] = 4; act_sel_in[1] = 1; act_sel_in[2] = 4; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 2; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 0; act_sel_in[14] = 1; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 4; act_sel_in[1] = 3; act_sel_in[2] = 1; act_sel_in[3] = 4; act_sel_in[4] = 0; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 1; act_sel_in[8] = 0; act_sel_in[9] = 4; act_sel_in[10] = 3; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 3; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=5; act_sel_in[0] = 4; act_sel_in[1] = 0; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 3; act_sel_in[5] = 0; act_sel_in[6] = 1; act_sel_in[7] = 3; act_sel_in[8] = 2; act_sel_in[9] = 1; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 2; act_sel_in[13] = 0; act_sel_in[14] = 1; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=4; act_sel_in[0] = 2; act_sel_in[1] = 2; act_sel_in[2] = 4; act_sel_in[3] = 2; act_sel_in[4] = 0; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 2; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 0; act_sel_in[11] = 3; act_sel_in[12] = 4; act_sel_in[13] = 3; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 0; act_sel_in[1] = 3; act_sel_in[2] = 1; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 2; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 2; act_sel_in[11] = 2; act_sel_in[12] = 4; act_sel_in[13] = 0; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=2; act_sel_in[0] = 3; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 3; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 0; act_sel_in[7] = 4; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 2; act_sel_in[12] = 4; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 3; act_sel_in[1] = 4; act_sel_in[2] = 1; act_sel_in[3] = 0; act_sel_in[4] = 0; act_sel_in[5] = 3; act_sel_in[6] = 0; act_sel_in[7] = 2; act_sel_in[8] = 2; act_sel_in[9] = 0; act_sel_in[10] = 3; act_sel_in[11] = 0; act_sel_in[12] = 3; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 4; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 4; act_sel_in[4] = 2; act_sel_in[5] = 2; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 0; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 


    #1 is_msb=1; column_idx=7; act[0] = -88; act[1] = -43; act[2] = -93; act[3] = -20; act[4] = 53; act[5] = 41; act[6] = 63; act[7] = -115; act[8] = 108; act[9] = 125; act[10] = 67; act[11] = 50; act[12] = -107; act[13] = -96; act[14] = -115; act[15] = 98; act[16] = -36; act[17] = -82; act[18] = -29; act[19] = 37; act[20] = -21; act[21] = -21; act[22] = -38; act[23] = -81; act[24] = 11; act[25] = -69; act[26] = -94; act[27] = 94; act[28] = 50; act[29] = -106; act[30] = -1; act[31] = 20; 
    act_sel_in[0] = 3; act_sel_in[1] = 0; act_sel_in[2] = 2; act_sel_in[3] = 2; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 2; act_sel_in[9] = 1; act_sel_in[10] = 3; act_sel_in[11] = 3; act_sel_in[12] = 0; act_sel_in[13] = 0; act_sel_in[14] = 1; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 3; act_sel_in[1] = 2; act_sel_in[2] = 2; act_sel_in[3] = 1; act_sel_in[4] = 0; act_sel_in[5] = 0; act_sel_in[6] = 4; act_sel_in[7] = 0; act_sel_in[8] = 3; act_sel_in[9] = 2; act_sel_in[10] = 1; act_sel_in[11] = 3; act_sel_in[12] = 3; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=5; act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 0; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 4; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 0; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 2; act_sel_in[12] = 3; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=4; act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 0; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 2; act_sel_in[7] = 3; act_sel_in[8] = 1; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 3; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 3; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=3; act_sel_in[0] = 1; act_sel_in[1] = 0; act_sel_in[2] = 1; act_sel_in[3] = 0; act_sel_in[4] = 4; act_sel_in[5] = 4; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 1; act_sel_in[9] = 1; act_sel_in[10] = 1; act_sel_in[11] = 0; act_sel_in[12] = 3; act_sel_in[13] = 3; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=2; act_sel_in[0] = 2; act_sel_in[1] = 4; act_sel_in[2] = 0; act_sel_in[3] = 3; act_sel_in[4] = 0; act_sel_in[5] = 3; act_sel_in[6] = 2; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 4; act_sel_in[10] = 4; act_sel_in[11] = 0; act_sel_in[12] = 4; act_sel_in[13] = 4; act_sel_in[14] = 1; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 3; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 3; act_sel_in[4] = 3; act_sel_in[5] = 4; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 2; act_sel_in[9] = 3; act_sel_in[10] = 3; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 1; act_sel_in[14] = 1; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=0; act_sel_in[0] = 4; act_sel_in[1] = 0; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 4; act_sel_in[9] = 2; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 3; act_sel_in[13] = 1; act_sel_in[14] = 3; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 


    #1 is_msb=1; column_idx=7; act[0] = 38; act[1] = 63; act[2] = 98; act[3] = -77; act[4] = 100; act[5] = 105; act[6] = -57; act[7] = -33; act[8] = -7; act[9] = 114; act[10] = -19; act[11] = -81; act[12] = 81; act[13] = 13; act[14] = 18; act[15] = 21; act[16] = -98; act[17] = 96; act[18] = -86; act[19] = -12; act[20] = 13; act[21] = 29; act[22] = -29; act[23] = 84; act[24] = 37; act[25] = -13; act[26] = -78; act[27] = -26; act[28] = 92; act[29] = 72; act[30] = 109; act[31] = -70; 
    act_sel_in[0] = 2; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 0; act_sel_in[4] = 2; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 4; act_sel_in[9] = 0; act_sel_in[10] = 4; act_sel_in[11] = 0; act_sel_in[12] = 3; act_sel_in[13] = 3; act_sel_in[14] = 3; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 4; act_sel_in[1] = 0; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 3; act_sel_in[5] = 4; act_sel_in[6] = 4; act_sel_in[7] = 4; act_sel_in[8] = 1; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 0; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=5; act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 4; act_sel_in[3] = 1; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 3; act_sel_in[11] = 0; act_sel_in[12] = 1; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=4; act_sel_in[0] = 0; act_sel_in[1] = 3; act_sel_in[2] = 4; act_sel_in[3] = 2; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 0; act_sel_in[7] = 1; act_sel_in[8] = 3; act_sel_in[9] = 1; act_sel_in[10] = 4; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 3; act_sel_in[14] = 1; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 0; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 0; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 2; act_sel_in[8] = 4; act_sel_in[9] = 3; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 1; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=2; act_sel_in[0] = 3; act_sel_in[1] = 4; act_sel_in[2] = 4; act_sel_in[3] = 0; act_sel_in[4] = 2; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 4; act_sel_in[8] = 1; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 4; act_sel_in[12] = 4; act_sel_in[13] = 0; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=1; act_sel_in[0] = 2; act_sel_in[1] = 3; act_sel_in[2] = 0; act_sel_in[3] = 3; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 4; act_sel_in[7] = 3; act_sel_in[8] = 1; act_sel_in[9] = 2; act_sel_in[10] = 0; act_sel_in[11] = 3; act_sel_in[12] = 2; act_sel_in[13] = 3; act_sel_in[14] = 4; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=0; act_sel_in[0] = 3; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 0; act_sel_in[4] = 0; act_sel_in[5] = 3; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 3; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 2; act_sel_in[12] = 3; act_sel_in[13] = 3; act_sel_in[14] = 1; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 


    #1 is_msb=1; column_idx=7; act[0] = 90; act[1] = -116; act[2] = 21; act[3] = 121; act[4] = -63; act[5] = 17; act[6] = -118; act[7] = -95; act[8] = -78; act[9] = -30; act[10] = 94; act[11] = 4; act[12] = -128; act[13] = 66; act[14] = -21; act[15] = 6; act[16] = -92; act[17] = 99; act[18] = -69; act[19] = 117; act[20] = -109; act[21] = 27; act[22] = 32; act[23] = 12; act[24] = 88; act[25] = -59; act[26] = 75; act[27] = 16; act[28] = 56; act[29] = 110; act[30] = -30; act[31] = 125; 
    act_sel_in[0] = 4; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 1; act_sel_in[4] = 3; act_sel_in[5] = 4; act_sel_in[6] = 4; act_sel_in[7] = 0; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 0; act_sel_in[11] = 2; act_sel_in[12] = 0; act_sel_in[13] = 0; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 0; act_sel_in[1] = 0; act_sel_in[2] = 2; act_sel_in[3] = 0; act_sel_in[4] = 0; act_sel_in[5] = 0; act_sel_in[6] = 4; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 1; act_sel_in[11] = 3; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 0; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=5; act_sel_in[0] = 0; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 2; act_sel_in[4] = 4; act_sel_in[5] = 1; act_sel_in[6] = 2; act_sel_in[7] = 4; act_sel_in[8] = 2; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 2; act_sel_in[14] = 1; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=4; act_sel_in[0] = 1; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 0; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 0; act_sel_in[10] = 0; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 0; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=3; act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 3; act_sel_in[5] = 1; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 4; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=2; act_sel_in[0] = 1; act_sel_in[1] = 4; act_sel_in[2] = 4; act_sel_in[3] = 3; act_sel_in[4] = 2; act_sel_in[5] = 4; act_sel_in[6] = 0; act_sel_in[7] = 2; act_sel_in[8] = 2; act_sel_in[9] = 3; act_sel_in[10] = 3; act_sel_in[11] = 3; act_sel_in[12] = 2; act_sel_in[13] = 3; act_sel_in[14] = 0; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 2; act_sel_in[1] = 4; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 4; act_sel_in[8] = 1; act_sel_in[9] = 2; act_sel_in[10] = 0; act_sel_in[11] = 2; act_sel_in[12] = 4; act_sel_in[13] = 4; act_sel_in[14] = 4; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 3; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 


    #1 is_msb=1; column_idx=7; act[0] = -35; act[1] = 87; act[2] = -112; act[3] = -69; act[4] = 51; act[5] = -46; act[6] = 25; act[7] = 79; act[8] = 51; act[9] = 19; act[10] = -17; act[11] = 105; act[12] = -58; act[13] = 55; act[14] = -120; act[15] = 98; act[16] = -109; act[17] = 34; act[18] = 40; act[19] = 108; act[20] = -128; act[21] = -114; act[22] = -119; act[23] = -23; act[24] = 11; act[25] = 78; act[26] = 55; act[27] = -106; act[28] = 61; act[29] = -123; act[30] = -125; act[31] = 70; 
    act_sel_in[0] = 1; act_sel_in[1] = 1; act_sel_in[2] = 0; act_sel_in[3] = 2; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 4; act_sel_in[8] = 4; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 1; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 3; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 2; act_sel_in[4] = 4; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 4; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 4; act_sel_in[14] = 1; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=5; act_sel_in[0] = 3; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 0; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 1; act_sel_in[10] = 4; act_sel_in[11] = 3; act_sel_in[12] = 3; act_sel_in[13] = 0; act_sel_in[14] = 1; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=4; act_sel_in[0] = 4; act_sel_in[1] = 4; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 3; act_sel_in[7] = 1; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 1; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=3; act_sel_in[0] = 1; act_sel_in[1] = 0; act_sel_in[2] = 1; act_sel_in[3] = 3; act_sel_in[4] = 2; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 2; act_sel_in[9] = 4; act_sel_in[10] = 4; act_sel_in[11] = 3; act_sel_in[12] = 1; act_sel_in[13] = 2; act_sel_in[14] = 3; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=2; act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 1; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 3; act_sel_in[1] = 1; act_sel_in[2] = 4; act_sel_in[3] = 1; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 0; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 1; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=0; act_sel_in[0] = 1; act_sel_in[1] = 0; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 2; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 3; act_sel_in[11] = 1; act_sel_in[12] = 0; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 


    #1 is_msb=1; column_idx=7; act[0] = 13; act[1] = 62; act[2] = -63; act[3] = -124; act[4] = 27; act[5] = -121; act[6] = -38; act[7] = -89; act[8] = -37; act[9] = -29; act[10] = 108; act[11] = -45; act[12] = 31; act[13] = 45; act[14] = -25; act[15] = 124; act[16] = 109; act[17] = -30; act[18] = 62; act[19] = -34; act[20] = 91; act[21] = 115; act[22] = -87; act[23] = -28; act[24] = -60; act[25] = -115; act[26] = 60; act[27] = -38; act[28] = -122; act[29] = -12; act[30] = 77; act[31] = 101; 
    act_sel_in[0] = 2; act_sel_in[1] = 4; act_sel_in[2] = 4; act_sel_in[3] = 2; act_sel_in[4] = 2; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 1; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 3; act_sel_in[9] = 4; act_sel_in[10] = 4; act_sel_in[11] = 4; act_sel_in[12] = 4; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=5; act_sel_in[0] = 3; act_sel_in[1] = 4; act_sel_in[2] = 1; act_sel_in[3] = 4; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 0; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 3; act_sel_in[12] = 4; act_sel_in[13] = 4; act_sel_in[14] = 3; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=4; act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 2; act_sel_in[3] = 3; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 1; act_sel_in[8] = 3; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 0; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 3; act_sel_in[1] = 3; act_sel_in[2] = 3; act_sel_in[3] = 4; act_sel_in[4] = 0; act_sel_in[5] = 4; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=2; act_sel_in[0] = 3; act_sel_in[1] = 4; act_sel_in[2] = 0; act_sel_in[3] = 2; act_sel_in[4] = 3; act_sel_in[5] = 4; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 3; act_sel_in[12] = 4; act_sel_in[13] = 4; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 2; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 0; act_sel_in[5] = 0; act_sel_in[6] = 1; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 2; act_sel_in[10] = 2; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 2; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 0; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 0; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 1; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 2; act_sel_in[10] = 0; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 


    #1 is_msb=1; column_idx=7; act[0] = -96; act[1] = -63; act[2] = 105; act[3] = -25; act[4] = -106; act[5] = -85; act[6] = 110; act[7] = 12; act[8] = -96; act[9] = 126; act[10] = 105; act[11] = -108; act[12] = -19; act[13] = 47; act[14] = -115; act[15] = 120; act[16] = 17; act[17] = -16; act[18] = 8; act[19] = 44; act[20] = 61; act[21] = 97; act[22] = 93; act[23] = -22; act[24] = 102; act[25] = 86; act[26] = 10; act[27] = 93; act[28] = 18; act[29] = -35; act[30] = 2; act[31] = -106; 
    act_sel_in[0] = 4; act_sel_in[1] = 3; act_sel_in[2] = 0; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 1; act_sel_in[11] = 1; act_sel_in[12] = 0; act_sel_in[13] = 0; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 2; act_sel_in[3] = 0; act_sel_in[4] = 0; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 4; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=5; act_sel_in[0] = 3; act_sel_in[1] = 3; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 3; act_sel_in[8] = 4; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 2; act_sel_in[14] = 1; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=4; act_sel_in[0] = 0; act_sel_in[1] = 3; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 1; act_sel_in[11] = 0; act_sel_in[12] = 4; act_sel_in[13] = 3; act_sel_in[14] = 1; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 4; act_sel_in[1] = 0; act_sel_in[2] = 3; act_sel_in[3] = 4; act_sel_in[4] = 0; act_sel_in[5] = 4; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 3; act_sel_in[11] = 3; act_sel_in[12] = 3; act_sel_in[13] = 2; act_sel_in[14] = 3; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=2; act_sel_in[0] = 4; act_sel_in[1] = 4; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 0; act_sel_in[7] = 4; act_sel_in[8] = 1; act_sel_in[9] = 0; act_sel_in[10] = 1; act_sel_in[11] = 3; act_sel_in[12] = 4; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 2; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 4; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 3; act_sel_in[11] = 2; act_sel_in[12] = 4; act_sel_in[13] = 3; act_sel_in[14] = 3; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 1; act_sel_in[4] = 3; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 2; act_sel_in[14] = 1; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 


    #1 is_msb=1; column_idx=7; act[0] = -50; act[1] = 59; act[2] = 4; act[3] = 6; act[4] = 10; act[5] = 6; act[6] = -100; act[7] = 29; act[8] = 22; act[9] = 20; act[10] = 3; act[11] = 57; act[12] = -23; act[13] = 87; act[14] = -81; act[15] = -81; act[16] = -27; act[17] = 97; act[18] = -59; act[19] = -29; act[20] = 99; act[21] = -21; act[22] = -37; act[23] = -4; act[24] = -92; act[25] = -77; act[26] = -77; act[27] = 74; act[28] = 113; act[29] = -23; act[30] = 62; act[31] = -82; 
    act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 1; act_sel_in[5] = 4; act_sel_in[6] = 3; act_sel_in[7] = 0; act_sel_in[8] = 2; act_sel_in[9] = 4; act_sel_in[10] = 3; act_sel_in[11] = 1; act_sel_in[12] = 0; act_sel_in[13] = 4; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 3; act_sel_in[1] = 0; act_sel_in[2] = 1; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 4; act_sel_in[8] = 4; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 0; act_sel_in[12] = 4; act_sel_in[13] = 3; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=5; act_sel_in[0] = 1; act_sel_in[1] = 4; act_sel_in[2] = 0; act_sel_in[3] = 2; act_sel_in[4] = 3; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 4; act_sel_in[9] = 3; act_sel_in[10] = 1; act_sel_in[11] = 3; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 4; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=4; act_sel_in[0] = 3; act_sel_in[1] = 0; act_sel_in[2] = 2; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 3; act_sel_in[8] = 4; act_sel_in[9] = 3; act_sel_in[10] = 4; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 0; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 3; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 3; act_sel_in[14] = 1; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=2; act_sel_in[0] = 3; act_sel_in[1] = 1; act_sel_in[2] = 2; act_sel_in[3] = 1; act_sel_in[4] = 3; act_sel_in[5] = 1; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 0; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 3; act_sel_in[12] = 2; act_sel_in[13] = 2; act_sel_in[14] = 1; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=1; act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 3; act_sel_in[5] = 4; act_sel_in[6] = 1; act_sel_in[7] = 4; act_sel_in[8] = 4; act_sel_in[9] = 2; act_sel_in[10] = 0; act_sel_in[11] = 4; act_sel_in[12] = 1; act_sel_in[13] = 3; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=0; act_sel_in[0] = 4; act_sel_in[1] = 1; act_sel_in[2] = 2; act_sel_in[3] = 1; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 0; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 3; act_sel_in[13] = 4; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 


    #1 is_msb=1; column_idx=7; act[0] = 72; act[1] = 57; act[2] = -121; act[3] = -111; act[4] = 1; act[5] = -44; act[6] = 51; act[7] = 72; act[8] = -105; act[9] = -60; act[10] = -56; act[11] = 95; act[12] = -99; act[13] = 81; act[14] = -66; act[15] = -47; act[16] = -102; act[17] = -12; act[18] = 26; act[19] = -80; act[20] = 11; act[21] = 52; act[22] = 73; act[23] = 127; act[24] = 84; act[25] = -97; act[26] = -84; act[27] = 50; act[28] = 90; act[29] = -1; act[30] = -126; act[31] = 50; 
    act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 2; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 0; act_sel_in[11] = 3; act_sel_in[12] = 1; act_sel_in[13] = 2; act_sel_in[14] = 0; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 2; act_sel_in[1] = 4; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 3; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 2; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 0; act_sel_in[14] = 3; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=5; act_sel_in[0] = 4; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 1; act_sel_in[4] = 0; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 1; act_sel_in[9] = 4; act_sel_in[10] = 3; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 0; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=4; act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 2; act_sel_in[3] = 2; act_sel_in[4] = 2; act_sel_in[5] = 4; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 2; act_sel_in[9] = 3; act_sel_in[10] = 4; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 0; act_sel_in[14] = 4; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 3; act_sel_in[1] = 1; act_sel_in[2] = 0; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 1; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 3; act_sel_in[13] = 4; act_sel_in[14] = 1; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=2; act_sel_in[0] = 2; act_sel_in[1] = 3; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 4; act_sel_in[9] = 2; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 4; act_sel_in[13] = 0; act_sel_in[14] = 0; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 2; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 3; act_sel_in[8] = 1; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 3; act_sel_in[14] = 0; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=0; act_sel_in[0] = 2; act_sel_in[1] = 0; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 2; act_sel_in[8] = 1; act_sel_in[9] = 4; act_sel_in[10] = 4; act_sel_in[11] = 2; act_sel_in[12] = 4; act_sel_in[13] = 1; act_sel_in[14] = 1; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 


    #1 is_msb=1; column_idx=7; act[0] = -82; act[1] = -113; act[2] = -72; act[3] = 86; act[4] = -89; act[5] = 70; act[6] = -65; act[7] = -3; act[8] = 9; act[9] = -120; act[10] = -101; act[11] = -60; act[12] = -17; act[13] = 52; act[14] = 124; act[15] = 61; act[16] = -47; act[17] = -31; act[18] = -76; act[19] = -58; act[20] = 49; act[21] = 66; act[22] = -66; act[23] = -68; act[24] = 18; act[25] = 42; act[26] = 116; act[27] = -125; act[28] = 72; act[29] = 51; act[30] = 99; act[31] = -114; 
    act_sel_in[0] = 3; act_sel_in[1] = 3; act_sel_in[2] = 1; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 4; act_sel_in[7] = 4; act_sel_in[8] = 2; act_sel_in[9] = 0; act_sel_in[10] = 2; act_sel_in[11] = 2; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 0; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 1; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 4; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 0; act_sel_in[14] = 2; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=5; act_sel_in[0] = 0; act_sel_in[1] = 3; act_sel_in[2] = 0; act_sel_in[3] = 0; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 1; act_sel_in[11] = 3; act_sel_in[12] = 2; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=4; act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 4; act_sel_in[3] = 4; act_sel_in[4] = 1; act_sel_in[5] = 4; act_sel_in[6] = 2; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=3; act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 2; act_sel_in[4] = 0; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 2; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 3; act_sel_in[12] = 1; act_sel_in[13] = 3; act_sel_in[14] = 4; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=2; act_sel_in[0] = 2; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 1; act_sel_in[4] = 3; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 3; act_sel_in[8] = 2; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 2; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 3; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 4; act_sel_in[4] = 0; act_sel_in[5] = 2; act_sel_in[6] = 0; act_sel_in[7] = 4; act_sel_in[8] = 1; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 3; act_sel_in[12] = 1; act_sel_in[13] = 4; act_sel_in[14] = 3; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 2; act_sel_in[1] = 3; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 3; act_sel_in[5] = 4; act_sel_in[6] = 1; act_sel_in[7] = 1; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 2; act_sel_in[11] = 3; act_sel_in[12] = 3; act_sel_in[13] = 4; act_sel_in[14] = 1; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 


    #1 is_msb=1; column_idx=7; act[0] = 50; act[1] = -51; act[2] = 32; act[3] = -41; act[4] = 33; act[5] = -77; act[6] = 22; act[7] = 61; act[8] = 60; act[9] = 4; act[10] = -106; act[11] = 2; act[12] = 54; act[13] = 12; act[14] = -113; act[15] = -43; act[16] = -72; act[17] = -10; act[18] = 44; act[19] = -44; act[20] = 99; act[21] = 96; act[22] = -115; act[23] = -102; act[24] = -20; act[25] = 8; act[26] = 114; act[27] = 44; act[28] = -20; act[29] = 8; act[30] = -100; act[31] = 56; 
    act_sel_in[0] = 4; act_sel_in[1] = 0; act_sel_in[2] = 4; act_sel_in[3] = 2; act_sel_in[4] = 2; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 2; act_sel_in[13] = 0; act_sel_in[14] = 0; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 0; act_sel_in[1] = 0; act_sel_in[2] = 0; act_sel_in[3] = 2; act_sel_in[4] = 0; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 3; act_sel_in[8] = 2; act_sel_in[9] = 3; act_sel_in[10] = 0; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 1; act_sel_in[14] = 0; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=5; act_sel_in[0] = 0; act_sel_in[1] = 1; act_sel_in[2] = 3; act_sel_in[3] = 2; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 0; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=4; act_sel_in[0] = 0; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 2; act_sel_in[4] = 2; act_sel_in[5] = 4; act_sel_in[6] = 3; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 4; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 3; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=3; act_sel_in[0] = 3; act_sel_in[1] = 2; act_sel_in[2] = 4; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 0; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 0; act_sel_in[11] = 0; act_sel_in[12] = 4; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=2; act_sel_in[0] = 4; act_sel_in[1] = 1; act_sel_in[2] = 0; act_sel_in[3] = 3; act_sel_in[4] = 2; act_sel_in[5] = 1; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 0; act_sel_in[10] = 4; act_sel_in[11] = 4; act_sel_in[12] = 3; act_sel_in[13] = 0; act_sel_in[14] = 3; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 1; act_sel_in[1] = 4; act_sel_in[2] = 0; act_sel_in[3] = 2; act_sel_in[4] = 0; act_sel_in[5] = 4; act_sel_in[6] = 2; act_sel_in[7] = 2; act_sel_in[8] = 2; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 1; act_sel_in[14] = 3; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 4; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 0; act_sel_in[4] = 0; act_sel_in[5] = 2; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 4; act_sel_in[10] = 0; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 3; act_sel_in[14] = 1; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 


    #1 is_msb=1; column_idx=7; act[0] = -119; act[1] = -31; act[2] = -64; act[3] = -110; act[4] = -79; act[5] = 34; act[6] = -128; act[7] = 59; act[8] = -84; act[9] = -109; act[10] = -48; act[11] = 85; act[12] = 17; act[13] = -55; act[14] = 27; act[15] = -16; act[16] = 53; act[17] = -64; act[18] = 85; act[19] = 91; act[20] = 101; act[21] = 29; act[22] = 35; act[23] = 121; act[24] = 67; act[25] = -11; act[26] = -54; act[27] = 15; act[28] = -86; act[29] = 57; act[30] = 29; act[31] = -120; 
    act_sel_in[0] = 3; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 0; act_sel_in[12] = 3; act_sel_in[13] = 3; act_sel_in[14] = 1; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 3; act_sel_in[1] = 2; act_sel_in[2] = 4; act_sel_in[3] = 3; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 0; act_sel_in[7] = 0; act_sel_in[8] = 4; act_sel_in[9] = 3; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=5; act_sel_in[0] = 2; act_sel_in[1] = 0; act_sel_in[2] = 1; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 0; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 2; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=4; act_sel_in[0] = 2; act_sel_in[1] = 4; act_sel_in[2] = 0; act_sel_in[3] = 3; act_sel_in[4] = 2; act_sel_in[5] = 3; act_sel_in[6] = 0; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 0; act_sel_in[10] = 3; act_sel_in[11] = 0; act_sel_in[12] = 3; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=3; act_sel_in[0] = 1; act_sel_in[1] = 1; act_sel_in[2] = 2; act_sel_in[3] = 0; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 4; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 2; act_sel_in[10] = 0; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=2; act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 1; act_sel_in[3] = 3; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 4; act_sel_in[7] = 4; act_sel_in[8] = 2; act_sel_in[9] = 3; act_sel_in[10] = 3; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 0; act_sel_in[14] = 1; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 4; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 4; act_sel_in[6] = 3; act_sel_in[7] = 0; act_sel_in[8] = 4; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 2; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 1; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=0; act_sel_in[0] = 3; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 3; act_sel_in[4] = 0; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 2; act_sel_in[8] = 3; act_sel_in[9] = 4; act_sel_in[10] = 0; act_sel_in[11] = 3; act_sel_in[12] = 4; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 


    #1 is_msb=1; column_idx=7; act[0] = 9; act[1] = -104; act[2] = 68; act[3] = 106; act[4] = -28; act[5] = -107; act[6] = -17; act[7] = 25; act[8] = -69; act[9] = 46; act[10] = 65; act[11] = 6; act[12] = 11; act[13] = 113; act[14] = 3; act[15] = 2; act[16] = -72; act[17] = -43; act[18] = -119; act[19] = -109; act[20] = -82; act[21] = -62; act[22] = -30; act[23] = -83; act[24] = 17; act[25] = 99; act[26] = 124; act[27] = 101; act[28] = 110; act[29] = -39; act[30] = 31; act[31] = 110; 
    act_sel_in[0] = 2; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 2; act_sel_in[5] = 4; act_sel_in[6] = 1; act_sel_in[7] = 1; act_sel_in[8] = 2; act_sel_in[9] = 1; act_sel_in[10] = 3; act_sel_in[11] = 3; act_sel_in[12] = 4; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 1; act_sel_in[1] = 1; act_sel_in[2] = 0; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 4; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=5; act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 2; act_sel_in[4] = 2; act_sel_in[5] = 3; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 2; act_sel_in[9] = 0; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 1; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=4; act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 4; act_sel_in[3] = 4; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 0; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 0; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 0; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 2; act_sel_in[1] = 0; act_sel_in[2] = 1; act_sel_in[3] = 0; act_sel_in[4] = 4; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 2; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 1; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 3; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=2; act_sel_in[0] = 0; act_sel_in[1] = 0; act_sel_in[2] = 0; act_sel_in[3] = 1; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 3; act_sel_in[12] = 3; act_sel_in[13] = 0; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 4; act_sel_in[8] = 4; act_sel_in[9] = 3; act_sel_in[10] = 4; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 3; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=0; act_sel_in[0] = 0; act_sel_in[1] = 0; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 2; act_sel_in[11] = 0; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 


    #1 is_msb=1; column_idx=7; act[0] = -41; act[1] = -99; act[2] = -76; act[3] = 64; act[4] = 100; act[5] = 116; act[6] = -88; act[7] = 14; act[8] = 115; act[9] = -36; act[10] = -3; act[11] = 1; act[12] = 102; act[13] = 49; act[14] = -42; act[15] = -90; act[16] = 38; act[17] = 64; act[18] = -113; act[19] = -105; act[20] = 20; act[21] = 94; act[22] = 22; act[23] = 17; act[24] = 85; act[25] = 50; act[26] = 127; act[27] = 6; act[28] = -113; act[29] = -20; act[30] = -103; act[31] = 39; 
    act_sel_in[0] = 1; act_sel_in[1] = 1; act_sel_in[2] = 4; act_sel_in[3] = 4; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 4; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 2; act_sel_in[11] = 2; act_sel_in[12] = 3; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 4; act_sel_in[1] = 4; act_sel_in[2] = 1; act_sel_in[3] = 3; act_sel_in[4] = 1; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 3; act_sel_in[9] = 1; act_sel_in[10] = 3; act_sel_in[11] = 3; act_sel_in[12] = 2; act_sel_in[13] = 0; act_sel_in[14] = 1; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=5; act_sel_in[0] = 0; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 3; act_sel_in[4] = 2; act_sel_in[5] = 3; act_sel_in[6] = 1; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 4; act_sel_in[10] = 0; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=4; act_sel_in[0] = 0; act_sel_in[1] = 1; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 2; act_sel_in[5] = 2; act_sel_in[6] = 0; act_sel_in[7] = 2; act_sel_in[8] = 2; act_sel_in[9] = 1; act_sel_in[10] = 4; act_sel_in[11] = 3; act_sel_in[12] = 3; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 0; act_sel_in[5] = 0; act_sel_in[6] = 0; act_sel_in[7] = 1; act_sel_in[8] = 1; act_sel_in[9] = 4; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 4; act_sel_in[14] = 2; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=2; act_sel_in[0] = 1; act_sel_in[1] = 1; act_sel_in[2] = 0; act_sel_in[3] = 1; act_sel_in[4] = 0; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 0; act_sel_in[10] = 2; act_sel_in[11] = 0; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 3; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=1; act_sel_in[0] = 0; act_sel_in[1] = 3; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 1; act_sel_in[7] = 1; act_sel_in[8] = 3; act_sel_in[9] = 2; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 0; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=0; act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 1; act_sel_in[3] = 4; act_sel_in[4] = 2; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 0; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 3; act_sel_in[11] = 3; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 4; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 


    #1 is_msb=1; column_idx=7; act[0] = -103; act[1] = 2; act[2] = 23; act[3] = -50; act[4] = 24; act[5] = 53; act[6] = 106; act[7] = -123; act[8] = 68; act[9] = -123; act[10] = 25; act[11] = 37; act[12] = 66; act[13] = 118; act[14] = -8; act[15] = 27; act[16] = 93; act[17] = -9; act[18] = 110; act[19] = -98; act[20] = -16; act[21] = -70; act[22] = 86; act[23] = 43; act[24] = -1; act[25] = -95; act[26] = 78; act[27] = 114; act[28] = 109; act[29] = 58; act[30] = -16; act[31] = 42; 
    act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 1; act_sel_in[4] = 1; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 1; act_sel_in[14] = 0; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 4; act_sel_in[6] = 3; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 2; act_sel_in[10] = 2; act_sel_in[11] = 4; act_sel_in[12] = 1; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=5; act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 4; act_sel_in[3] = 4; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 3; act_sel_in[9] = 0; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 1; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=4; act_sel_in[0] = 4; act_sel_in[1] = 0; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 2; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 4; act_sel_in[9] = 0; act_sel_in[10] = 4; act_sel_in[11] = 3; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 4; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 4; act_sel_in[9] = 0; act_sel_in[10] = 4; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 3; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=2; act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 2; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 4; act_sel_in[8] = 4; act_sel_in[9] = 4; act_sel_in[10] = 0; act_sel_in[11] = 4; act_sel_in[12] = 3; act_sel_in[13] = 4; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=1; act_sel_in[0] = 3; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 3; act_sel_in[4] = 0; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 2; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 2; act_sel_in[14] = 3; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 3; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 1; act_sel_in[8] = 1; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 


    #1 is_msb=1; column_idx=7; act[0] = -32; act[1] = -71; act[2] = 9; act[3] = 125; act[4] = -42; act[5] = -68; act[6] = 26; act[7] = -126; act[8] = 100; act[9] = 56; act[10] = 72; act[11] = 94; act[12] = 89; act[13] = -100; act[14] = 1; act[15] = -6; act[16] = 89; act[17] = -47; act[18] = -40; act[19] = 75; act[20] = 28; act[21] = 33; act[22] = -91; act[23] = 57; act[24] = 19; act[25] = 2; act[26] = -78; act[27] = -67; act[28] = -11; act[29] = 91; act[30] = 110; act[31] = -53; 
    act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 4; act_sel_in[6] = 0; act_sel_in[7] = 0; act_sel_in[8] = 4; act_sel_in[9] = 0; act_sel_in[10] = 3; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 4; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 4; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 2; act_sel_in[10] = 3; act_sel_in[11] = 3; act_sel_in[12] = 1; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=5; act_sel_in[0] = 1; act_sel_in[1] = 4; act_sel_in[2] = 4; act_sel_in[3] = 0; act_sel_in[4] = 2; act_sel_in[5] = 1; act_sel_in[6] = 0; act_sel_in[7] = 2; act_sel_in[8] = 3; act_sel_in[9] = 0; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 0; act_sel_in[13] = 4; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=4; act_sel_in[0] = 0; act_sel_in[1] = 0; act_sel_in[2] = 2; act_sel_in[3] = 2; act_sel_in[4] = 2; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 2; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 4; act_sel_in[12] = 1; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=3; act_sel_in[0] = 3; act_sel_in[1] = 1; act_sel_in[2] = 4; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 0; act_sel_in[6] = 0; act_sel_in[7] = 1; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 2; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 1; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=2; act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 1; act_sel_in[9] = 3; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 1; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=1; act_sel_in[0] = 3; act_sel_in[1] = 1; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 3; act_sel_in[5] = 1; act_sel_in[6] = 2; act_sel_in[7] = 4; act_sel_in[8] = 2; act_sel_in[9] = 0; act_sel_in[10] = 4; act_sel_in[11] = 4; act_sel_in[12] = 1; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=0; act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 1; act_sel_in[3] = 3; act_sel_in[4] = 4; act_sel_in[5] = 1; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 2; act_sel_in[9] = 0; act_sel_in[10] = 2; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 2; act_sel_in[14] = 1; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 


    #1 is_msb=1; column_idx=7; act[0] = 89; act[1] = 47; act[2] = -33; act[3] = -45; act[4] = 36; act[5] = 101; act[6] = -108; act[7] = -63; act[8] = 80; act[9] = -62; act[10] = 107; act[11] = 116; act[12] = 39; act[13] = -11; act[14] = -15; act[15] = 46; act[16] = -61; act[17] = 71; act[18] = -43; act[19] = -82; act[20] = 113; act[21] = -11; act[22] = 93; act[23] = -118; act[24] = -47; act[25] = -18; act[26] = 100; act[27] = 59; act[28] = 112; act[29] = 35; act[30] = -83; act[31] = -116; 
    act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 1; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 1; act_sel_in[8] = 4; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 0; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 3; act_sel_in[1] = 2; act_sel_in[2] = 2; act_sel_in[3] = 1; act_sel_in[4] = 3; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 3; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 1; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=5; act_sel_in[0] = 1; act_sel_in[1] = 1; act_sel_in[2] = 2; act_sel_in[3] = 1; act_sel_in[4] = 0; act_sel_in[5] = 1; act_sel_in[6] = 3; act_sel_in[7] = 0; act_sel_in[8] = 3; act_sel_in[9] = 0; act_sel_in[10] = 4; act_sel_in[11] = 4; act_sel_in[12] = 3; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=4; act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 4; act_sel_in[3] = 1; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 4; act_sel_in[7] = 0; act_sel_in[8] = 3; act_sel_in[9] = 2; act_sel_in[10] = 1; act_sel_in[11] = 4; act_sel_in[12] = 3; act_sel_in[13] = 0; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 2; act_sel_in[1] = 0; act_sel_in[2] = 2; act_sel_in[3] = 3; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 2; act_sel_in[7] = 3; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 3; act_sel_in[11] = 2; act_sel_in[12] = 0; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=2; act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 2; act_sel_in[3] = 2; act_sel_in[4] = 0; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 0; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 3; act_sel_in[14] = 1; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=1; act_sel_in[0] = 3; act_sel_in[1] = 4; act_sel_in[2] = 0; act_sel_in[3] = 2; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 0; act_sel_in[8] = 4; act_sel_in[9] = 2; act_sel_in[10] = 3; act_sel_in[11] = 1; act_sel_in[12] = 0; act_sel_in[13] = 2; act_sel_in[14] = 1; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 4; act_sel_in[3] = 3; act_sel_in[4] = 4; act_sel_in[5] = 4; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 2; act_sel_in[9] = 0; act_sel_in[10] = 3; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 1; act_sel_in[14] = 0; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 


    #1 is_msb=1; column_idx=7; act[0] = 14; act[1] = -50; act[2] = 14; act[3] = 36; act[4] = 95; act[5] = 62; act[6] = 24; act[7] = 22; act[8] = -59; act[9] = -26; act[10] = 30; act[11] = -49; act[12] = 33; act[13] = -126; act[14] = 91; act[15] = -53; act[16] = 85; act[17] = 17; act[18] = 102; act[19] = 4; act[20] = -25; act[21] = -44; act[22] = -12; act[23] = -117; act[24] = -53; act[25] = -101; act[26] = -52; act[27] = 24; act[28] = -4; act[29] = 26; act[30] = 54; act[31] = -29; 
    act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 3; act_sel_in[7] = 1; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 3; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 0; act_sel_in[1] = 0; act_sel_in[2] = 2; act_sel_in[3] = 0; act_sel_in[4] = 0; act_sel_in[5] = 0; act_sel_in[6] = 0; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 1; act_sel_in[12] = 2; act_sel_in[13] = 0; act_sel_in[14] = 0; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=5; act_sel_in[0] = 3; act_sel_in[1] = 3; act_sel_in[2] = 4; act_sel_in[3] = 4; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 0; act_sel_in[7] = 1; act_sel_in[8] = 1; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 4; act_sel_in[14] = 3; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=4; act_sel_in[0] = 3; act_sel_in[1] = 0; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 1; act_sel_in[9] = 2; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 4; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 0; act_sel_in[5] = 4; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 2; act_sel_in[9] = 1; act_sel_in[10] = 3; act_sel_in[11] = 3; act_sel_in[12] = 0; act_sel_in[13] = 4; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=2; act_sel_in[0] = 1; act_sel_in[1] = 0; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=1; act_sel_in[0] = 4; act_sel_in[1] = 3; act_sel_in[2] = 4; act_sel_in[3] = 0; act_sel_in[4] = 0; act_sel_in[5] = 4; act_sel_in[6] = 0; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 3; act_sel_in[11] = 1; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 4; act_sel_in[8] = 2; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 3; act_sel_in[12] = 2; act_sel_in[13] = 1; act_sel_in[14] = 1; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 


    #1 is_msb=1; column_idx=7; act[0] = 5; act[1] = -108; act[2] = 0; act[3] = -60; act[4] = 60; act[5] = 37; act[6] = 103; act[7] = 44; act[8] = 6; act[9] = -118; act[10] = 28; act[11] = 101; act[12] = 36; act[13] = -31; act[14] = -109; act[15] = 20; act[16] = -87; act[17] = 94; act[18] = -23; act[19] = 39; act[20] = 6; act[21] = 38; act[22] = 52; act[23] = 117; act[24] = 95; act[25] = 53; act[26] = 96; act[27] = 103; act[28] = 101; act[29] = -124; act[30] = -22; act[31] = 12; 
    act_sel_in[0] = 2; act_sel_in[1] = 2; act_sel_in[2] = 2; act_sel_in[3] = 2; act_sel_in[4] = 3; act_sel_in[5] = 1; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 3; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 1; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 1; act_sel_in[1] = 4; act_sel_in[2] = 1; act_sel_in[3] = 3; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=5; act_sel_in[0] = 4; act_sel_in[1] = 4; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 2; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 3; act_sel_in[9] = 0; act_sel_in[10] = 3; act_sel_in[11] = 0; act_sel_in[12] = 1; act_sel_in[13] = 3; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=4; act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 4; act_sel_in[3] = 4; act_sel_in[4] = 1; act_sel_in[5] = 4; act_sel_in[6] = 2; act_sel_in[7] = 2; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=3; act_sel_in[0] = 4; act_sel_in[1] = 1; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 1; act_sel_in[5] = 4; act_sel_in[6] = 3; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 3; act_sel_in[11] = 3; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=2; act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 1; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=1; act_sel_in[0] = 0; act_sel_in[1] = 1; act_sel_in[2] = 3; act_sel_in[3] = 4; act_sel_in[4] = 1; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 2; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 3; act_sel_in[11] = 1; act_sel_in[12] = 0; act_sel_in[13] = 4; act_sel_in[14] = 2; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 3; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 2; act_sel_in[6] = 3; act_sel_in[7] = 1; act_sel_in[8] = 2; act_sel_in[9] = 0; act_sel_in[10] = 3; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 1; act_sel_in[14] = 1; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 


    #1 is_msb=1; column_idx=7; act[0] = -8; act[1] = 120; act[2] = -39; act[3] = -77; act[4] = 29; act[5] = -20; act[6] = -1; act[7] = -69; act[8] = -109; act[9] = 35; act[10] = -69; act[11] = -94; act[12] = 18; act[13] = 28; act[14] = 46; act[15] = 64; act[16] = -116; act[17] = 18; act[18] = -121; act[19] = 14; act[20] = 7; act[21] = -127; act[22] = -13; act[23] = 127; act[24] = 29; act[25] = -77; act[26] = 95; act[27] = -17; act[28] = -50; act[29] = 1; act[30] = -2; act[31] = -53; 
    act_sel_in[0] = 0; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 3; act_sel_in[4] = 2; act_sel_in[5] = 0; act_sel_in[6] = 1; act_sel_in[7] = 3; act_sel_in[8] = 2; act_sel_in[9] = 3; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 3; act_sel_in[13] = 3; act_sel_in[14] = 3; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 2; act_sel_in[1] = 4; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 0; act_sel_in[5] = 0; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 4; act_sel_in[10] = 4; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 1; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=5; act_sel_in[0] = 2; act_sel_in[1] = 0; act_sel_in[2] = 3; act_sel_in[3] = 4; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 2; act_sel_in[11] = 0; act_sel_in[12] = 3; act_sel_in[13] = 0; act_sel_in[14] = 3; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=4; act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 3; act_sel_in[9] = 4; act_sel_in[10] = 3; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=3; act_sel_in[0] = 3; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 3; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 4; act_sel_in[7] = 4; act_sel_in[8] = 2; act_sel_in[9] = 0; act_sel_in[10] = 0; act_sel_in[11] = 3; act_sel_in[12] = 3; act_sel_in[13] = 1; act_sel_in[14] = 0; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=2; act_sel_in[0] = 1; act_sel_in[1] = 4; act_sel_in[2] = 0; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 0; act_sel_in[7] = 1; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 3; act_sel_in[11] = 1; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 2; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=1; act_sel_in[0] = 1; act_sel_in[1] = 1; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 4; act_sel_in[8] = 4; act_sel_in[9] = 3; act_sel_in[10] = 3; act_sel_in[11] = 3; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 2; act_sel_in[4] = 0; act_sel_in[5] = 1; act_sel_in[6] = 3; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 4; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 


    #1 is_msb=1; column_idx=7; act[0] = 25; act[1] = -123; act[2] = -101; act[3] = -92; act[4] = -25; act[5] = -95; act[6] = -74; act[7] = 52; act[8] = -33; act[9] = 121; act[10] = -6; act[11] = -85; act[12] = 90; act[13] = -17; act[14] = 59; act[15] = 97; act[16] = 66; act[17] = -20; act[18] = -71; act[19] = -102; act[20] = -24; act[21] = 60; act[22] = 102; act[23] = -105; act[24] = 43; act[25] = 70; act[26] = -88; act[27] = 18; act[28] = 50; act[29] = -29; act[30] = 96; act[31] = -18; 
    act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 0; act_sel_in[5] = 0; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 1; act_sel_in[9] = 4; act_sel_in[10] = 3; act_sel_in[11] = 0; act_sel_in[12] = 1; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 3; act_sel_in[1] = 3; act_sel_in[2] = 4; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 4; act_sel_in[11] = 3; act_sel_in[12] = 4; act_sel_in[13] = 1; act_sel_in[14] = 3; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=5; act_sel_in[0] = 4; act_sel_in[1] = 1; act_sel_in[2] = 2; act_sel_in[3] = 0; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 0; act_sel_in[7] = 1; act_sel_in[8] = 1; act_sel_in[9] = 2; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 2; act_sel_in[13] = 2; act_sel_in[14] = 3; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=4; act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 0; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 0; act_sel_in[7] = 4; act_sel_in[8] = 2; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 2; act_sel_in[14] = 1; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 0; act_sel_in[1] = 1; act_sel_in[2] = 4; act_sel_in[3] = 2; act_sel_in[4] = 2; act_sel_in[5] = 0; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 2; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 1; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=2; act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 4; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 1; act_sel_in[9] = 0; act_sel_in[10] = 3; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 0; act_sel_in[14] = 1; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 3; act_sel_in[1] = 2; act_sel_in[2] = 1; act_sel_in[3] = 3; act_sel_in[4] = 2; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 4; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 4; act_sel_in[12] = 1; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 3; act_sel_in[1] = 1; act_sel_in[2] = 0; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 1; act_sel_in[6] = 0; act_sel_in[7] = 1; act_sel_in[8] = 1; act_sel_in[9] = 4; act_sel_in[10] = 3; act_sel_in[11] = 2; act_sel_in[12] = 4; act_sel_in[13] = 0; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 


    #1 is_msb=1; column_idx=7; act[0] = 38; act[1] = -68; act[2] = -114; act[3] = 92; act[4] = 110; act[5] = 121; act[6] = -1; act[7] = -126; act[8] = 24; act[9] = 40; act[10] = 16; act[11] = -81; act[12] = -91; act[13] = -58; act[14] = -123; act[15] = 29; act[16] = -42; act[17] = -38; act[18] = 75; act[19] = 58; act[20] = -110; act[21] = -104; act[22] = -25; act[23] = 0; act[24] = 50; act[25] = 37; act[26] = -66; act[27] = 101; act[28] = -73; act[29] = -123; act[30] = 39; act[31] = -30; 
    act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 0; act_sel_in[4] = 2; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 4; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 1; act_sel_in[1] = 0; act_sel_in[2] = 1; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 1; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 0; act_sel_in[10] = 4; act_sel_in[11] = 0; act_sel_in[12] = 3; act_sel_in[13] = 1; act_sel_in[14] = 1; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=5; act_sel_in[0] = 2; act_sel_in[1] = 2; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 3; act_sel_in[9] = 4; act_sel_in[10] = 4; act_sel_in[11] = 0; act_sel_in[12] = 1; act_sel_in[13] = 0; act_sel_in[14] = 1; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=4; act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 1; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 1; act_sel_in[6] = 1; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 4; act_sel_in[12] = 4; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=3; act_sel_in[0] = 0; act_sel_in[1] = 0; act_sel_in[2] = 4; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 0; act_sel_in[9] = 2; act_sel_in[10] = 3; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 1; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=2; act_sel_in[0] = 0; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 2; act_sel_in[9] = 0; act_sel_in[10] = 0; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 3; act_sel_in[14] = 1; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=1; act_sel_in[0] = 2; act_sel_in[1] = 3; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 4; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 3; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 2; act_sel_in[9] = 3; act_sel_in[10] = 1; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 2; act_sel_in[14] = 1; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 


    #1 is_msb=1; column_idx=7; act[0] = 117; act[1] = -90; act[2] = 3; act[3] = 105; act[4] = 23; act[5] = -26; act[6] = -40; act[7] = 6; act[8] = -27; act[9] = 112; act[10] = -86; act[11] = 108; act[12] = -84; act[13] = -110; act[14] = -30; act[15] = -49; act[16] = -92; act[17] = -41; act[18] = 123; act[19] = -32; act[20] = -108; act[21] = 14; act[22] = -21; act[23] = -43; act[24] = 58; act[25] = 92; act[26] = -30; act[27] = -104; act[28] = -29; act[29] = -109; act[30] = 116; act[31] = -68; 
    act_sel_in[0] = 4; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 0; act_sel_in[7] = 4; act_sel_in[8] = 1; act_sel_in[9] = 1; act_sel_in[10] = 3; act_sel_in[11] = 0; act_sel_in[12] = 4; act_sel_in[13] = 1; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 4; act_sel_in[1] = 1; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 0; act_sel_in[9] = 2; act_sel_in[10] = 1; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 0; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=5; act_sel_in[0] = 2; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 2; act_sel_in[8] = 1; act_sel_in[9] = 1; act_sel_in[10] = 1; act_sel_in[11] = 3; act_sel_in[12] = 3; act_sel_in[13] = 0; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=4; act_sel_in[0] = 0; act_sel_in[1] = 3; act_sel_in[2] = 4; act_sel_in[3] = 4; act_sel_in[4] = 0; act_sel_in[5] = 3; act_sel_in[6] = 4; act_sel_in[7] = 0; act_sel_in[8] = 3; act_sel_in[9] = 2; act_sel_in[10] = 1; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 1; act_sel_in[10] = 3; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 3; act_sel_in[14] = 1; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=2; act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 2; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 3; act_sel_in[8] = 1; act_sel_in[9] = 2; act_sel_in[10] = 3; act_sel_in[11] = 3; act_sel_in[12] = 1; act_sel_in[13] = 3; act_sel_in[14] = 1; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=1; act_sel_in[0] = 0; act_sel_in[1] = 0; act_sel_in[2] = 2; act_sel_in[3] = 0; act_sel_in[4] = 2; act_sel_in[5] = 2; act_sel_in[6] = 0; act_sel_in[7] = 2; act_sel_in[8] = 3; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 0; act_sel_in[12] = 1; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 1; act_sel_in[1] = 4; act_sel_in[2] = 0; act_sel_in[3] = 2; act_sel_in[4] = 3; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 1; act_sel_in[8] = 2; act_sel_in[9] = 0; act_sel_in[10] = 0; act_sel_in[11] = 3; act_sel_in[12] = 4; act_sel_in[13] = 0; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 


    #1 is_msb=1; column_idx=7; act[0] = -59; act[1] = -80; act[2] = 12; act[3] = -14; act[4] = -104; act[5] = 102; act[6] = 21; act[7] = -62; act[8] = 61; act[9] = 115; act[10] = 25; act[11] = -71; act[12] = -35; act[13] = 17; act[14] = 118; act[15] = -103; act[16] = -69; act[17] = -44; act[18] = -15; act[19] = -118; act[20] = -21; act[21] = -70; act[22] = -113; act[23] = 78; act[24] = -1; act[25] = 14; act[26] = 9; act[27] = -74; act[28] = 90; act[29] = 122; act[30] = -61; act[31] = -12; 
    act_sel_in[0] = 4; act_sel_in[1] = 1; act_sel_in[2] = 2; act_sel_in[3] = 3; act_sel_in[4] = 2; act_sel_in[5] = 1; act_sel_in[6] = 0; act_sel_in[7] = 1; act_sel_in[8] = 1; act_sel_in[9] = 2; act_sel_in[10] = 0; act_sel_in[11] = 0; act_sel_in[12] = 4; act_sel_in[13] = 1; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 2; act_sel_in[1] = 0; act_sel_in[2] = 0; act_sel_in[3] = 0; act_sel_in[4] = 2; act_sel_in[5] = 1; act_sel_in[6] = 2; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 0; act_sel_in[14] = 0; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=5; act_sel_in[0] = 3; act_sel_in[1] = 4; act_sel_in[2] = 0; act_sel_in[3] = 2; act_sel_in[4] = 3; act_sel_in[5] = 1; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 3; act_sel_in[12] = 1; act_sel_in[13] = 1; act_sel_in[14] = 1; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=4; act_sel_in[0] = 1; act_sel_in[1] = 0; act_sel_in[2] = 1; act_sel_in[3] = 3; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 3; act_sel_in[11] = 2; act_sel_in[12] = 4; act_sel_in[13] = 4; act_sel_in[14] = 3; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 2; act_sel_in[1] = 0; act_sel_in[2] = 4; act_sel_in[3] = 0; act_sel_in[4] = 2; act_sel_in[5] = 3; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 2; act_sel_in[9] = 0; act_sel_in[10] = 1; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 0; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=2; act_sel_in[0] = 3; act_sel_in[1] = 1; act_sel_in[2] = 4; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 4; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 3; act_sel_in[12] = 2; act_sel_in[13] = 0; act_sel_in[14] = 2; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 3; act_sel_in[1] = 0; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 2; act_sel_in[9] = 0; act_sel_in[10] = 0; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 0; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=0; act_sel_in[0] = 3; act_sel_in[1] = 1; act_sel_in[2] = 4; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 2; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 


    #1 is_msb=1; column_idx=7; act[0] = -127; act[1] = 106; act[2] = 116; act[3] = 47; act[4] = 106; act[5] = -108; act[6] = -86; act[7] = -84; act[8] = 53; act[9] = -87; act[10] = 70; act[11] = 25; act[12] = -44; act[13] = 50; act[14] = 4; act[15] = -125; act[16] = -11; act[17] = -87; act[18] = -100; act[19] = 101; act[20] = -25; act[21] = -77; act[22] = -54; act[23] = -126; act[24] = 37; act[25] = -49; act[26] = 123; act[27] = 80; act[28] = 80; act[29] = -106; act[30] = -76; act[31] = -112; 
    act_sel_in[0] = 4; act_sel_in[1] = 3; act_sel_in[2] = 1; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 0; act_sel_in[6] = 1; act_sel_in[7] = 1; act_sel_in[8] = 3; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 4; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 3; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 0; act_sel_in[5] = 3; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 2; act_sel_in[9] = 4; act_sel_in[10] = 4; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=5; act_sel_in[0] = 3; act_sel_in[1] = 0; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 3; act_sel_in[9] = 0; act_sel_in[10] = 0; act_sel_in[11] = 0; act_sel_in[12] = 3; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=4; act_sel_in[0] = 4; act_sel_in[1] = 4; act_sel_in[2] = 0; act_sel_in[3] = 2; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 4; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=3; act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 4; act_sel_in[6] = 0; act_sel_in[7] = 1; act_sel_in[8] = 3; act_sel_in[9] = 2; act_sel_in[10] = 3; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 0; act_sel_in[14] = 3; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=2; act_sel_in[0] = 4; act_sel_in[1] = 0; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 3; act_sel_in[5] = 4; act_sel_in[6] = 2; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 0; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 1; act_sel_in[5] = 0; act_sel_in[6] = 0; act_sel_in[7] = 2; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 4; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 0; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=0; act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 4; act_sel_in[6] = 0; act_sel_in[7] = 0; act_sel_in[8] = 4; act_sel_in[9] = 2; act_sel_in[10] = 1; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 


    #1 is_msb=1; column_idx=7; act[0] = -29; act[1] = -125; act[2] = 28; act[3] = -33; act[4] = -115; act[5] = 88; act[6] = -2; act[7] = 56; act[8] = -77; act[9] = -96; act[10] = 84; act[11] = 54; act[12] = 88; act[13] = 37; act[14] = -96; act[15] = -25; act[16] = -127; act[17] = -71; act[18] = 121; act[19] = -64; act[20] = 28; act[21] = -45; act[22] = -51; act[23] = 85; act[24] = 126; act[25] = 89; act[26] = 79; act[27] = -83; act[28] = 104; act[29] = -118; act[30] = -84; act[31] = -30; 
    act_sel_in[0] = 2; act_sel_in[1] = 4; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 0; act_sel_in[5] = 3; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 0; act_sel_in[10] = 3; act_sel_in[11] = 1; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 1; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 3; act_sel_in[1] = 0; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 3; act_sel_in[5] = 0; act_sel_in[6] = 1; act_sel_in[7] = 1; act_sel_in[8] = 4; act_sel_in[9] = 0; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 4; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=5; act_sel_in[0] = 4; act_sel_in[1] = 1; act_sel_in[2] = 2; act_sel_in[3] = 2; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 4; act_sel_in[9] = 4; act_sel_in[10] = 0; act_sel_in[11] = 3; act_sel_in[12] = 3; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=4; act_sel_in[0] = 0; act_sel_in[1] = 0; act_sel_in[2] = 4; act_sel_in[3] = 4; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 0; act_sel_in[7] = 0; act_sel_in[8] = 4; act_sel_in[9] = 0; act_sel_in[10] = 0; act_sel_in[11] = 3; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 3; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=3; act_sel_in[0] = 2; act_sel_in[1] = 2; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 4; act_sel_in[5] = 4; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 2; act_sel_in[10] = 0; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 3; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=2; act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 4; act_sel_in[10] = 4; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 0; act_sel_in[14] = 2; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 4; act_sel_in[1] = 1; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 1; act_sel_in[7] = 4; act_sel_in[8] = 4; act_sel_in[9] = 3; act_sel_in[10] = 3; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=0; act_sel_in[0] = 1; act_sel_in[1] = 1; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 0; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 1; act_sel_in[8] = 1; act_sel_in[9] = 2; act_sel_in[10] = 0; act_sel_in[11] = 4; act_sel_in[12] = 4; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 


    #1 is_msb=1; column_idx=7; act[0] = 20; act[1] = -73; act[2] = -50; act[3] = 27; act[4] = 86; act[5] = 84; act[6] = 28; act[7] = -31; act[8] = 73; act[9] = -103; act[10] = 42; act[11] = -67; act[12] = 40; act[13] = 86; act[14] = 11; act[15] = 21; act[16] = -119; act[17] = -10; act[18] = 104; act[19] = -47; act[20] = 100; act[21] = 114; act[22] = 12; act[23] = -5; act[24] = 73; act[25] = -19; act[26] = 96; act[27] = -106; act[28] = -49; act[29] = -8; act[30] = -94; act[31] = 66; 
    act_sel_in[0] = 3; act_sel_in[1] = 3; act_sel_in[2] = 4; act_sel_in[3] = 3; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 3; act_sel_in[9] = 0; act_sel_in[10] = 0; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 1; act_sel_in[1] = 0; act_sel_in[2] = 2; act_sel_in[3] = 3; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 2; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 4; act_sel_in[14] = 4; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=5; act_sel_in[0] = 1; act_sel_in[1] = 1; act_sel_in[2] = 4; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 1; act_sel_in[6] = 1; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 4; act_sel_in[11] = 2; act_sel_in[12] = 3; act_sel_in[13] = 1; act_sel_in[14] = 3; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=4; act_sel_in[0] = 0; act_sel_in[1] = 1; act_sel_in[2] = 0; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 0; act_sel_in[7] = 0; act_sel_in[8] = 3; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 2; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=3; act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 3; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 4; act_sel_in[8] = 2; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 3; act_sel_in[12] = 1; act_sel_in[13] = 3; act_sel_in[14] = 4; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=2; act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 4; act_sel_in[3] = 1; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 0; act_sel_in[7] = 1; act_sel_in[8] = 3; act_sel_in[9] = 1; act_sel_in[10] = 3; act_sel_in[11] = 0; act_sel_in[12] = 3; act_sel_in[13] = 2; act_sel_in[14] = 1; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 3; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 1; act_sel_in[9] = 3; act_sel_in[10] = 1; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 0; act_sel_in[14] = 3; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 0; act_sel_in[5] = 3; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 1; act_sel_in[9] = 1; act_sel_in[10] = 3; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 4; act_sel_in[14] = 2; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 


    #1 is_msb=1; column_idx=7; act[0] = 26; act[1] = -11; act[2] = 127; act[3] = 17; act[4] = -88; act[5] = -82; act[6] = -107; act[7] = 101; act[8] = -39; act[9] = -89; act[10] = -80; act[11] = 21; act[12] = -68; act[13] = 4; act[14] = -98; act[15] = -12; act[16] = -16; act[17] = -75; act[18] = 124; act[19] = -6; act[20] = 55; act[21] = 79; act[22] = -52; act[23] = 74; act[24] = -37; act[25] = 95; act[26] = 60; act[27] = -114; act[28] = 30; act[29] = 92; act[30] = 120; act[31] = 74; 
    act_sel_in[0] = 3; act_sel_in[1] = 0; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 1; act_sel_in[7] = 3; act_sel_in[8] = 1; act_sel_in[9] = 0; act_sel_in[10] = 0; act_sel_in[11] = 3; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 4; act_sel_in[1] = 4; act_sel_in[2] = 1; act_sel_in[3] = 3; act_sel_in[4] = 0; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 2; act_sel_in[11] = 4; act_sel_in[12] = 4; act_sel_in[13] = 1; act_sel_in[14] = 1; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=5; act_sel_in[0] = 1; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 2; act_sel_in[10] = 3; act_sel_in[11] = 2; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 3; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=4; act_sel_in[0] = 2; act_sel_in[1] = 2; act_sel_in[2] = 2; act_sel_in[3] = 1; act_sel_in[4] = 3; act_sel_in[5] = 4; act_sel_in[6] = 1; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 4; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 0; act_sel_in[14] = 1; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 1; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 3; act_sel_in[11] = 4; act_sel_in[12] = 4; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=2; act_sel_in[0] = 4; act_sel_in[1] = 0; act_sel_in[2] = 0; act_sel_in[3] = 2; act_sel_in[4] = 0; act_sel_in[5] = 2; act_sel_in[6] = 3; act_sel_in[7] = 1; act_sel_in[8] = 4; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 3; act_sel_in[14] = 1; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=1; act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 4; act_sel_in[3] = 3; act_sel_in[4] = 0; act_sel_in[5] = 1; act_sel_in[6] = 2; act_sel_in[7] = 3; act_sel_in[8] = 3; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 2; act_sel_in[12] = 4; act_sel_in[13] = 4; act_sel_in[14] = 1; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 2; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 2; act_sel_in[4] = 2; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 3; act_sel_in[8] = 4; act_sel_in[9] = 4; act_sel_in[10] = 0; act_sel_in[11] = 3; act_sel_in[12] = 3; act_sel_in[13] = 4; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 





    #15 $stop;
  end

  always #1 clk = ~clk;

endmodule

`endif