`ifndef __vert_32_tb_V__
`define __vert_32_tb_V__

`include "mac_unit_Vert_32_no_mul.v"

module vert_32_tb;
    
    parameter DATA_WIDTH    = 8;
    parameter VEC_LENGTH    = 32;
    parameter MUX_SEL_WIDTH = 3;
    parameter SUM_ACT_WIDTH = $clog2(VEC_LENGTH) + DATA_WIDTH - 2;
    parameter ACC_WIDTH     = DATA_WIDTH + 16;
    parameter RESULT_WIDTH  = 2*DATA_WIDTH;

    logic                               clk;
    logic                               reset;
    logic                               en_acc;
    logic                               load_accum;

    logic signed   [DATA_WIDTH-1:0]     act         [VEC_LENGTH-1:0];   // input activation (signed)
    logic          [MUX_SEL_WIDTH-1:0]  act_sel_in  [VEC_LENGTH/2-1:0]; // input activation MUX select signal
    logic                               act_val_in  [VEC_LENGTH/2-1:0]; // whether activation is valid
    logic signed   [SUM_ACT_WIDTH-1:0]  sum_act  [VEC_LENGTH/8-1:0]; // sum of a group of activations (signed)

    logic          [2:0]                column_idx;    // current column index for shifting 
    logic                               is_msb;        // specify if the current column is MSB
    logic                               is_skip_zero [VEC_LENGTH/8-1:0];  // specify if skip bit 0
    
    logic signed   [ACC_WIDTH-1:0]      accum_prev;
    logic signed   [RESULT_WIDTH-1:0]   result;

    mac_unit_Vert_32_no_mul_clk #(DATA_WIDTH, VEC_LENGTH, MUX_SEL_WIDTH, SUM_ACT_WIDTH, ACC_WIDTH) dut (.*);

  initial
    $monitor ("out=%b", result);

  initial begin
    `ifdef SIMULATE 
      $vcdpluson;
      $vcdplusmemon;
    `endif

    #0 clk = 0; reset = 1;  en_acc = 0;
    #1 reset = 0; en_acc = 1; load_accum = 0; accum_prev = 0; sum_act[1]=100; sum_act[2]=100; sum_act[3]=100; sum_act[4]=100;

    #1.25 is_msb_in=1; column_idx_in=7; act[0] = 10; act[1] = 83; act[2] = -24; act[3] = 103; act[4] = 47; act[5] = -93; act[6] = -99; act[7] = -88; act[8] = 98; act[9] = 93; act[10] = 108; act[11] = -3; act[12] = 33; act[13] = 61; act[14] = -71; act[15] = -30; act[16] = 5; act[17] = -18; act[18] = 118; act[19] = 39; act[20] = 36; act[21] = 108; act[22] = 36; act[23] = 59; act[24] = -1; act[25] = 74; act[26] = 24; act[27] = -101; act[28] = 108; act[29] = -12; act[30] = -117; act[31] = -56; 
act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 1; act_sel_in[3] = 3; act_sel_in[4] = 0; act_sel_in[5] = 2; act_sel_in[6] = 0; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 0; act_sel_in[12] = 4; act_sel_in[13] = 3; act_sel_in[14] = 4; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 is_msb_in=0; column_idx_in=6; act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 2; act_sel_in[3] = 1; act_sel_in[4] = 0; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 2; act_sel_in[13] = 0; act_sel_in[14] = 0; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=5; act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 0; act_sel_in[3] = 1; act_sel_in[4] = 0; act_sel_in[5] = 2; act_sel_in[6] = 3; act_sel_in[7] = 2; act_sel_in[8] = 4; act_sel_in[9] = 2; act_sel_in[10] = 3; act_sel_in[11] = 2; act_sel_in[12] = 0; act_sel_in[13] = 0; act_sel_in[14] = 1; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=4; act_sel_in[0] = 4; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 0; act_sel_in[4] = 2; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 3; act_sel_in[8] = 2; act_sel_in[9] = 3; act_sel_in[10] = 2; act_sel_in[11] = 2; act_sel_in[12] = 4; act_sel_in[13] = 1; act_sel_in[14] = 1; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=3; act_sel_in[0] = 3; act_sel_in[1] = 3; act_sel_in[2] = 0; act_sel_in[3] = 3; act_sel_in[4] = 0; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 4; act_sel_in[10] = 3; act_sel_in[11] = 2; act_sel_in[12] = 0; act_sel_in[13] = 2; act_sel_in[14] = 3; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=2; act_sel_in[0] = 3; act_sel_in[1] = 4; act_sel_in[2] = 0; act_sel_in[3] = 2; act_sel_in[4] = 4; act_sel_in[5] = 1; act_sel_in[6] = 0; act_sel_in[7] = 1; act_sel_in[8] = 1; act_sel_in[9] = 3; act_sel_in[10] = 0; act_sel_in[11] = 4; act_sel_in[12] = 1; act_sel_in[13] = 1; act_sel_in[14] = 3; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=1; act_sel_in[0] = 4; act_sel_in[1] = 0; act_sel_in[2] = 3; act_sel_in[3] = 2; act_sel_in[4] = 2; act_sel_in[5] = 3; act_sel_in[6] = 0; act_sel_in[7] = 2; act_sel_in[8] = 2; act_sel_in[9] = 1; act_sel_in[10] = 1; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 3; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=0; act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 4; act_sel_in[3] = 1; act_sel_in[4] = 0; act_sel_in[5] = 0; act_sel_in[6] = 0; act_sel_in[7] = 3; act_sel_in[8] = 1; act_sel_in[9] = 3; act_sel_in[10] = 4; act_sel_in[11] = 0; act_sel_in[12] = 1; act_sel_in[13] = 0; act_sel_in[14] = 3; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 


#1.25 is_msb_in=1; column_idx_in=7; act[0] = 103; act[1] = 53; act[2] = 64; act[3] = 55; act[4] = -81; act[5] = -72; act[6] = -101; act[7] = 44; act[8] = 107; act[9] = 113; act[10] = -45; act[11] = 82; act[12] = 86; act[13] = 5; act[14] = -3; act[15] = -100; act[16] = -45; act[17] = -77; act[18] = -90; act[19] = -105; act[20] = -17; act[21] = 66; act[22] = -124; act[23] = 103; act[24] = -58; act[25] = -89; act[26] = 41; act[27] = -47; act[28] = -23; act[29] = -52; act[30] = -59; act[31] = -27; 
act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 1; act_sel_in[4] = 1; act_sel_in[5] = 4; act_sel_in[6] = 0; act_sel_in[7] = 4; act_sel_in[8] = 2; act_sel_in[9] = 1; act_sel_in[10] = 1; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 2; act_sel_in[14] = 1; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 is_msb_in=0; column_idx_in=6; act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 1; act_sel_in[3] = 3; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 0; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 3; act_sel_in[12] = 2; act_sel_in[13] = 2; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=5; act_sel_in[0] = 3; act_sel_in[1] = 3; act_sel_in[2] = 3; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 2; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 4; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 4; act_sel_in[14] = 3; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=4; act_sel_in[0] = 2; act_sel_in[1] = 2; act_sel_in[2] = 2; act_sel_in[3] = 0; act_sel_in[4] = 0; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 2; act_sel_in[9] = 3; act_sel_in[10] = 0; act_sel_in[11] = 0; act_sel_in[12] = 1; act_sel_in[13] = 4; act_sel_in[14] = 1; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=3; act_sel_in[0] = 0; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 0; act_sel_in[4] = 0; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 3; act_sel_in[9] = 2; act_sel_in[10] = 2; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=2; act_sel_in[0] = 4; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 3; act_sel_in[4] = 2; act_sel_in[5] = 4; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 3; act_sel_in[9] = 0; act_sel_in[10] = 3; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 3; act_sel_in[14] = 1; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=1; act_sel_in[0] = 4; act_sel_in[1] = 1; act_sel_in[2] = 2; act_sel_in[3] = 3; act_sel_in[4] = 3; act_sel_in[5] = 1; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 1; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 4; act_sel_in[14] = 1; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=0; act_sel_in[0] = 0; act_sel_in[1] = 1; act_sel_in[2] = 2; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 4; act_sel_in[6] = 1; act_sel_in[7] = 3; act_sel_in[8] = 3; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 2; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 


#1.25 is_msb_in=1; column_idx_in=7; act[0] = -87; act[1] = -14; act[2] = 20; act[3] = 111; act[4] = 0; act[5] = -97; act[6] = -84; act[7] = 15; act[8] = -107; act[9] = 97; act[10] = 14; act[11] = -9; act[12] = 116; act[13] = 17; act[14] = -114; act[15] = 117; act[16] = -24; act[17] = 46; act[18] = -19; act[19] = -107; act[20] = 79; act[21] = 26; act[22] = 43; act[23] = 98; act[24] = -3; act[25] = 98; act[26] = -123; act[27] = 105; act[28] = -18; act[29] = 30; act[30] = -19; act[31] = -106; 
act_sel_in[0] = 2; act_sel_in[1] = 0; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 3; act_sel_in[12] = 0; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 is_msb_in=0; column_idx_in=6; act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 4; act_sel_in[6] = 0; act_sel_in[7] = 1; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 3; act_sel_in[11] = 4; act_sel_in[12] = 3; act_sel_in[13] = 0; act_sel_in[14] = 0; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=5; act_sel_in[0] = 2; act_sel_in[1] = 2; act_sel_in[2] = 2; act_sel_in[3] = 1; act_sel_in[4] = 0; act_sel_in[5] = 1; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 3; act_sel_in[12] = 3; act_sel_in[13] = 0; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=4; act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 1; act_sel_in[6] = 2; act_sel_in[7] = 2; act_sel_in[8] = 1; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 1; act_sel_in[12] = 0; act_sel_in[13] = 4; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=3; act_sel_in[0] = 4; act_sel_in[1] = 4; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 2; act_sel_in[5] = 0; act_sel_in[6] = 4; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 0; act_sel_in[10] = 0; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 0; act_sel_in[14] = 1; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=2; act_sel_in[0] = 2; act_sel_in[1] = 4; act_sel_in[2] = 0; act_sel_in[3] = 3; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 0; act_sel_in[7] = 0; act_sel_in[8] = 4; act_sel_in[9] = 0; act_sel_in[10] = 1; act_sel_in[11] = 4; act_sel_in[12] = 4; act_sel_in[13] = 3; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=1; act_sel_in[0] = 0; act_sel_in[1] = 3; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 0; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 1; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=0; act_sel_in[0] = 3; act_sel_in[1] = 0; act_sel_in[2] = 1; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 4; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 4; act_sel_in[9] = 0; act_sel_in[10] = 3; act_sel_in[11] = 3; act_sel_in[12] = 0; act_sel_in[13] = 0; act_sel_in[14] = 0; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 


#1.25 is_msb_in=1; column_idx_in=7; act[0] = 111; act[1] = -24; act[2] = 30; act[3] = 77; act[4] = -98; act[5] = 20; act[6] = 26; act[7] = -91; act[8] = -94; act[9] = 74; act[10] = -65; act[11] = 33; act[12] = -35; act[13] = 94; act[14] = -18; act[15] = -68; act[16] = 72; act[17] = -32; act[18] = 84; act[19] = 60; act[20] = -88; act[21] = -68; act[22] = 66; act[23] = -5; act[24] = -30; act[25] = -123; act[26] = 81; act[27] = -36; act[28] = -72; act[29] = 85; act[30] = -127; act[31] = 54; 
act_sel_in[0] = 4; act_sel_in[1] = 0; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 0; act_sel_in[11] = 3; act_sel_in[12] = 3; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 is_msb_in=0; column_idx_in=6; act_sel_in[0] = 2; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 0; act_sel_in[11] = 4; act_sel_in[12] = 3; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=5; act_sel_in[0] = 2; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 0; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 1; act_sel_in[11] = 0; act_sel_in[12] = 3; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=4; act_sel_in[0] = 3; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 1; act_sel_in[7] = 1; act_sel_in[8] = 2; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 1; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=3; act_sel_in[0] = 0; act_sel_in[1] = 3; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 2; act_sel_in[5] = 3; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 1; act_sel_in[11] = 0; act_sel_in[12] = 1; act_sel_in[13] = 4; act_sel_in[14] = 4; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=2; act_sel_in[0] = 3; act_sel_in[1] = 4; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 1; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=1; act_sel_in[0] = 4; act_sel_in[1] = 1; act_sel_in[2] = 0; act_sel_in[3] = 3; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 3; act_sel_in[11] = 2; act_sel_in[12] = 3; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=0; act_sel_in[0] = 0; act_sel_in[1] = 0; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 3; act_sel_in[11] = 1; act_sel_in[12] = 2; act_sel_in[13] = 3; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 


#1.25 is_msb_in=1; column_idx_in=7; act[0] = 109; act[1] = -89; act[2] = 125; act[3] = -96; act[4] = -39; act[5] = 78; act[6] = -81; act[7] = 120; act[8] = -80; act[9] = 17; act[10] = -10; act[11] = 7; act[12] = -13; act[13] = -13; act[14] = -75; act[15] = -31; act[16] = -128; act[17] = -106; act[18] = -27; act[19] = -48; act[20] = 35; act[21] = 119; act[22] = 34; act[23] = 44; act[24] = -39; act[25] = 62; act[26] = 95; act[27] = 26; act[28] = -57; act[29] = -103; act[30] = -23; act[31] = -61; 
act_sel_in[0] = 0; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 3; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 2; act_sel_in[7] = 2; act_sel_in[8] = 0; act_sel_in[9] = 2; act_sel_in[10] = 2; act_sel_in[11] = 3; act_sel_in[12] = 2; act_sel_in[13] = 0; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 is_msb_in=0; column_idx_in=6; act_sel_in[0] = 1; act_sel_in[1] = 0; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 2; act_sel_in[7] = 4; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 2; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=5; act_sel_in[0] = 1; act_sel_in[1] = 4; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 2; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 2; act_sel_in[8] = 2; act_sel_in[9] = 0; act_sel_in[10] = 1; act_sel_in[11] = 1; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=4; act_sel_in[0] = 3; act_sel_in[1] = 3; act_sel_in[2] = 1; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 1; act_sel_in[8] = 1; act_sel_in[9] = 3; act_sel_in[10] = 0; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 0; act_sel_in[14] = 3; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=3; act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 4; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 2; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 4; act_sel_in[12] = 4; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=2; act_sel_in[0] = 3; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 4; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 4; act_sel_in[10] = 0; act_sel_in[11] = 2; act_sel_in[12] = 3; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=1; act_sel_in[0] = 1; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 3; act_sel_in[4] = 2; act_sel_in[5] = 3; act_sel_in[6] = 4; act_sel_in[7] = 4; act_sel_in[8] = 1; act_sel_in[9] = 3; act_sel_in[10] = 3; act_sel_in[11] = 0; act_sel_in[12] = 3; act_sel_in[13] = 1; act_sel_in[14] = 1; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=0; act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 0; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 1; act_sel_in[9] = 2; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 


#1.25 is_msb_in=1; column_idx_in=7; act[0] = 44; act[1] = 71; act[2] = -124; act[3] = 73; act[4] = -126; act[5] = 75; act[6] = 38; act[7] = 22; act[8] = -13; act[9] = -30; act[10] = -10; act[11] = 75; act[12] = 84; act[13] = 68; act[14] = 8; act[15] = -78; act[16] = -31; act[17] = 10; act[18] = 127; act[19] = -88; act[20] = 28; act[21] = 44; act[22] = 72; act[23] = 121; act[24] = 96; act[25] = -70; act[26] = 56; act[27] = 52; act[28] = 31; act[29] = -107; act[30] = 109; act[31] = -52; 
act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 0; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 0; act_sel_in[7] = 1; act_sel_in[8] = 4; act_sel_in[9] = 3; act_sel_in[10] = 1; act_sel_in[11] = 3; act_sel_in[12] = 1; act_sel_in[13] = 0; act_sel_in[14] = 3; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 is_msb_in=0; column_idx_in=6; act_sel_in[0] = 2; act_sel_in[1] = 3; act_sel_in[2] = 0; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 0; act_sel_in[6] = 4; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 3; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 3; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=5; act_sel_in[0] = 1; act_sel_in[1] = 1; act_sel_in[2] = 0; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 3; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 1; act_sel_in[9] = 0; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 4; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=4; act_sel_in[0] = 1; act_sel_in[1] = 0; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 4; act_sel_in[6] = 0; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 3; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 4; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=3; act_sel_in[0] = 3; act_sel_in[1] = 0; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 1; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 2; act_sel_in[9] = 4; act_sel_in[10] = 0; act_sel_in[11] = 3; act_sel_in[12] = 4; act_sel_in[13] = 3; act_sel_in[14] = 1; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=2; act_sel_in[0] = 3; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 0; act_sel_in[5] = 4; act_sel_in[6] = 4; act_sel_in[7] = 0; act_sel_in[8] = 4; act_sel_in[9] = 0; act_sel_in[10] = 3; act_sel_in[11] = 0; act_sel_in[12] = 1; act_sel_in[13] = 4; act_sel_in[14] = 1; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=1; act_sel_in[0] = 4; act_sel_in[1] = 0; act_sel_in[2] = 4; act_sel_in[3] = 4; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 2; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 3; act_sel_in[14] = 1; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=0; act_sel_in[0] = 4; act_sel_in[1] = 0; act_sel_in[2] = 1; act_sel_in[3] = 3; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 4; act_sel_in[8] = 4; act_sel_in[9] = 2; act_sel_in[10] = 1; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 3; act_sel_in[14] = 3; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 


#1.25 is_msb_in=1; column_idx_in=7; act[0] = 94; act[1] = 61; act[2] = -124; act[3] = -118; act[4] = 125; act[5] = -81; act[6] = 84; act[7] = -18; act[8] = -11; act[9] = 56; act[10] = -9; act[11] = 41; act[12] = 32; act[13] = 111; act[14] = 109; act[15] = 99; act[16] = 110; act[17] = -128; act[18] = -55; act[19] = -68; act[20] = 120; act[21] = 7; act[22] = -74; act[23] = -99; act[24] = 100; act[25] = -87; act[26] = 9; act[27] = -41; act[28] = 33; act[29] = -28; act[30] = 8; act[31] = 6; 
act_sel_in[0] = 1; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 3; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 3; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 3; act_sel_in[11] = 3; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 is_msb_in=0; column_idx_in=6; act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 3; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 0; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=5; act_sel_in[0] = 2; act_sel_in[1] = 0; act_sel_in[2] = 0; act_sel_in[3] = 2; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 3; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=4; act_sel_in[0] = 4; act_sel_in[1] = 0; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 1; act_sel_in[5] = 0; act_sel_in[6] = 4; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 2; act_sel_in[11] = 0; act_sel_in[12] = 3; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=3; act_sel_in[0] = 4; act_sel_in[1] = 1; act_sel_in[2] = 3; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 3; act_sel_in[8] = 4; act_sel_in[9] = 4; act_sel_in[10] = 3; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 0; act_sel_in[14] = 2; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=2; act_sel_in[0] = 3; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 2; act_sel_in[5] = 1; act_sel_in[6] = 2; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 1; act_sel_in[10] = 3; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 0; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=1; act_sel_in[0] = 3; act_sel_in[1] = 3; act_sel_in[2] = 0; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 4; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 4; act_sel_in[9] = 0; act_sel_in[10] = 1; act_sel_in[11] = 3; act_sel_in[12] = 1; act_sel_in[13] = 4; act_sel_in[14] = 3; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=0; act_sel_in[0] = 4; act_sel_in[1] = 3; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 4; act_sel_in[6] = 3; act_sel_in[7] = 0; act_sel_in[8] = 4; act_sel_in[9] = 2; act_sel_in[10] = 3; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 3; act_sel_in[14] = 1; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 


#1.25 is_msb_in=1; column_idx_in=7; act[0] = 80; act[1] = 24; act[2] = -99; act[3] = 67; act[4] = 95; act[5] = 73; act[6] = 100; act[7] = -58; act[8] = 41; act[9] = 33; act[10] = -66; act[11] = 109; act[12] = -89; act[13] = 18; act[14] = -107; act[15] = -23; act[16] = 37; act[17] = -88; act[18] = -124; act[19] = -77; act[20] = -79; act[21] = -85; act[22] = 32; act[23] = -66; act[24] = -107; act[25] = 14; act[26] = 93; act[27] = -106; act[28] = -116; act[29] = -38; act[30] = -25; act[31] = -32; 
act_sel_in[0] = 3; act_sel_in[1] = 4; act_sel_in[2] = 4; act_sel_in[3] = 4; act_sel_in[4] = 3; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 4; act_sel_in[9] = 3; act_sel_in[10] = 4; act_sel_in[11] = 3; act_sel_in[12] = 3; act_sel_in[13] = 0; act_sel_in[14] = 4; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 is_msb_in=0; column_idx_in=6; act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 0; act_sel_in[3] = 2; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 1; act_sel_in[7] = 3; act_sel_in[8] = 3; act_sel_in[9] = 0; act_sel_in[10] = 4; act_sel_in[11] = 0; act_sel_in[12] = 1; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=5; act_sel_in[0] = 3; act_sel_in[1] = 2; act_sel_in[2] = 4; act_sel_in[3] = 0; act_sel_in[4] = 4; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 2; act_sel_in[10] = 0; act_sel_in[11] = 0; act_sel_in[12] = 1; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=4; act_sel_in[0] = 3; act_sel_in[1] = 0; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 1; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 4; act_sel_in[10] = 0; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 0; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=3; act_sel_in[0] = 2; act_sel_in[1] = 2; act_sel_in[2] = 2; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 0; act_sel_in[8] = 4; act_sel_in[9] = 0; act_sel_in[10] = 1; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 1; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=2; act_sel_in[0] = 2; act_sel_in[1] = 0; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 1; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 2; act_sel_in[10] = 0; act_sel_in[11] = 2; act_sel_in[12] = 4; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=1; act_sel_in[0] = 3; act_sel_in[1] = 2; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 0; act_sel_in[5] = 1; act_sel_in[6] = 3; act_sel_in[7] = 2; act_sel_in[8] = 4; act_sel_in[9] = 4; act_sel_in[10] = 3; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=0; act_sel_in[0] = 4; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 2; act_sel_in[4] = 0; act_sel_in[5] = 4; act_sel_in[6] = 0; act_sel_in[7] = 2; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 3; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 2; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 


#1.25 is_msb_in=1; column_idx_in=7; act[0] = 75; act[1] = 30; act[2] = -63; act[3] = 35; act[4] = 106; act[5] = 33; act[6] = 17; act[7] = -5; act[8] = -8; act[9] = -66; act[10] = -67; act[11] = 112; act[12] = -89; act[13] = 78; act[14] = 83; act[15] = 12; act[16] = -57; act[17] = 25; act[18] = -46; act[19] = -60; act[20] = 91; act[21] = 59; act[22] = 75; act[23] = 11; act[24] = -38; act[25] = -51; act[26] = -74; act[27] = 60; act[28] = 121; act[29] = -106; act[30] = -49; act[31] = -52; 
act_sel_in[0] = 2; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 2; act_sel_in[7] = 3; act_sel_in[8] = 3; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 3; act_sel_in[12] = 3; act_sel_in[13] = 0; act_sel_in[14] = 3; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 is_msb_in=0; column_idx_in=6; act_sel_in[0] = 2; act_sel_in[1] = 4; act_sel_in[2] = 1; act_sel_in[3] = 0; act_sel_in[4] = 4; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 2; act_sel_in[11] = 3; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 3; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=5; act_sel_in[0] = 3; act_sel_in[1] = 3; act_sel_in[2] = 1; act_sel_in[3] = 0; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 2; act_sel_in[7] = 4; act_sel_in[8] = 1; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 0; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=4; act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 3; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 4; act_sel_in[10] = 3; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 2; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=3; act_sel_in[0] = 0; act_sel_in[1] = 1; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 0; act_sel_in[7] = 1; act_sel_in[8] = 3; act_sel_in[9] = 2; act_sel_in[10] = 2; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=2; act_sel_in[0] = 4; act_sel_in[1] = 3; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 3; act_sel_in[8] = 1; act_sel_in[9] = 4; act_sel_in[10] = 4; act_sel_in[11] = 2; act_sel_in[12] = 4; act_sel_in[13] = 3; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=1; act_sel_in[0] = 4; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 2; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 1; act_sel_in[9] = 3; act_sel_in[10] = 0; act_sel_in[11] = 3; act_sel_in[12] = 0; act_sel_in[13] = 0; act_sel_in[14] = 4; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=0; act_sel_in[0] = 2; act_sel_in[1] = 3; act_sel_in[2] = 1; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 4; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 3; act_sel_in[9] = 0; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 0; act_sel_in[14] = 3; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 


#1.25 is_msb_in=1; column_idx_in=7; act[0] = -112; act[1] = -78; act[2] = -10; act[3] = 67; act[4] = -5; act[5] = 42; act[6] = -70; act[7] = 117; act[8] = -79; act[9] = -59; act[10] = -35; act[11] = 32; act[12] = 120; act[13] = 104; act[14] = 110; act[15] = -44; act[16] = -31; act[17] = -72; act[18] = 83; act[19] = -116; act[20] = 41; act[21] = -59; act[22] = 17; act[23] = 35; act[24] = 58; act[25] = 80; act[26] = -46; act[27] = 15; act[28] = 76; act[29] = -21; act[30] = 6; act[31] = 49; 
act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 1; act_sel_in[8] = 4; act_sel_in[9] = 0; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 0; act_sel_in[13] = 4; act_sel_in[14] = 1; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 is_msb_in=0; column_idx_in=6; act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 1; act_sel_in[7] = 3; act_sel_in[8] = 2; act_sel_in[9] = 0; act_sel_in[10] = 2; act_sel_in[11] = 4; act_sel_in[12] = 3; act_sel_in[13] = 4; act_sel_in[14] = 2; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=5; act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 1; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 0; act_sel_in[7] = 1; act_sel_in[8] = 4; act_sel_in[9] = 0; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=4; act_sel_in[0] = 0; act_sel_in[1] = 3; act_sel_in[2] = 0; act_sel_in[3] = 2; act_sel_in[4] = 3; act_sel_in[5] = 0; act_sel_in[6] = 0; act_sel_in[7] = 3; act_sel_in[8] = 2; act_sel_in[9] = 3; act_sel_in[10] = 0; act_sel_in[11] = 3; act_sel_in[12] = 2; act_sel_in[13] = 3; act_sel_in[14] = 3; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=3; act_sel_in[0] = 4; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 0; act_sel_in[4] = 2; act_sel_in[5] = 4; act_sel_in[6] = 4; act_sel_in[7] = 4; act_sel_in[8] = 1; act_sel_in[9] = 3; act_sel_in[10] = 0; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=2; act_sel_in[0] = 4; act_sel_in[1] = 3; act_sel_in[2] = 3; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 2; act_sel_in[9] = 3; act_sel_in[10] = 2; act_sel_in[11] = 4; act_sel_in[12] = 1; act_sel_in[13] = 2; act_sel_in[14] = 0; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=1; act_sel_in[0] = 4; act_sel_in[1] = 1; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 4; act_sel_in[8] = 2; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 2; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=0; act_sel_in[0] = 1; act_sel_in[1] = 1; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 3; act_sel_in[5] = 4; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 1; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 3; act_sel_in[14] = 1; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 


#1.25 is_msb_in=1; column_idx_in=7; act[0] = -22; act[1] = -82; act[2] = -54; act[3] = -99; act[4] = 21; act[5] = -99; act[6] = -121; act[7] = -31; act[8] = 8; act[9] = -119; act[10] = -16; act[11] = 117; act[12] = 19; act[13] = 103; act[14] = -60; act[15] = -67; act[16] = 96; act[17] = 121; act[18] = -122; act[19] = 61; act[20] = 40; act[21] = -63; act[22] = 95; act[23] = -74; act[24] = -27; act[25] = 43; act[26] = 70; act[27] = 127; act[28] = -64; act[29] = 25; act[30] = 101; act[31] = -77; 
act_sel_in[0] = 0; act_sel_in[1] = 1; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 0; act_sel_in[5] = 1; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 2; act_sel_in[9] = 3; act_sel_in[10] = 1; act_sel_in[11] = 4; act_sel_in[12] = 4; act_sel_in[13] = 1; act_sel_in[14] = 1; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 is_msb_in=0; column_idx_in=6; act_sel_in[0] = 4; act_sel_in[1] = 1; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 3; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 3; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 3; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 0; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=5; act_sel_in[0] = 2; act_sel_in[1] = 2; act_sel_in[2] = 4; act_sel_in[3] = 2; act_sel_in[4] = 2; act_sel_in[5] = 4; act_sel_in[6] = 4; act_sel_in[7] = 0; act_sel_in[8] = 3; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=4; act_sel_in[0] = 4; act_sel_in[1] = 3; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 0; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 2; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 2; act_sel_in[14] = 3; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=3; act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 2; act_sel_in[8] = 4; act_sel_in[9] = 4; act_sel_in[10] = 3; act_sel_in[11] = 3; act_sel_in[12] = 3; act_sel_in[13] = 4; act_sel_in[14] = 1; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=2; act_sel_in[0] = 2; act_sel_in[1] = 3; act_sel_in[2] = 0; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 3; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 3; act_sel_in[9] = 1; act_sel_in[10] = 1; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 1; act_sel_in[14] = 1; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=1; act_sel_in[0] = 3; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 3; act_sel_in[9] = 2; act_sel_in[10] = 3; act_sel_in[11] = 3; act_sel_in[12] = 1; act_sel_in[13] = 3; act_sel_in[14] = 3; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=0; act_sel_in[0] = 0; act_sel_in[1] = 1; act_sel_in[2] = 3; act_sel_in[3] = 4; act_sel_in[4] = 0; act_sel_in[5] = 4; act_sel_in[6] = 3; act_sel_in[7] = 0; act_sel_in[8] = 3; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 


#1.25 is_msb_in=1; column_idx_in=7; act[0] = 91; act[1] = 48; act[2] = 112; act[3] = 26; act[4] = 35; act[5] = -104; act[6] = 122; act[7] = 116; act[8] = -46; act[9] = 56; act[10] = -12; act[11] = 53; act[12] = -49; act[13] = 53; act[14] = -100; act[15] = 112; act[16] = -38; act[17] = -37; act[18] = -37; act[19] = 109; act[20] = 103; act[21] = 115; act[22] = 81; act[23] = -90; act[24] = 35; act[25] = -36; act[26] = -32; act[27] = -109; act[28] = -111; act[29] = 15; act[30] = 58; act[31] = 34; 
act_sel_in[0] = 4; act_sel_in[1] = 3; act_sel_in[2] = 4; act_sel_in[3] = 2; act_sel_in[4] = 0; act_sel_in[5] = 1; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 2; act_sel_in[11] = 3; act_sel_in[12] = 3; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 is_msb_in=0; column_idx_in=6; act_sel_in[0] = 4; act_sel_in[1] = 3; act_sel_in[2] = 4; act_sel_in[3] = 0; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 1; act_sel_in[11] = 4; act_sel_in[12] = 3; act_sel_in[13] = 0; act_sel_in[14] = 3; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=5; act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 1; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 1; act_sel_in[9] = 0; act_sel_in[10] = 2; act_sel_in[11] = 3; act_sel_in[12] = 3; act_sel_in[13] = 0; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=4; act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 0; act_sel_in[3] = 3; act_sel_in[4] = 3; act_sel_in[5] = 4; act_sel_in[6] = 2; act_sel_in[7] = 2; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 2; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 0; act_sel_in[14] = 2; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=3; act_sel_in[0] = 0; act_sel_in[1] = 3; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 1; act_sel_in[6] = 1; act_sel_in[7] = 3; act_sel_in[8] = 4; act_sel_in[9] = 2; act_sel_in[10] = 3; act_sel_in[11] = 1; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 1; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=2; act_sel_in[0] = 3; act_sel_in[1] = 1; act_sel_in[2] = 0; act_sel_in[3] = 0; act_sel_in[4] = 4; act_sel_in[5] = 1; act_sel_in[6] = 2; act_sel_in[7] = 3; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 4; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=1; act_sel_in[0] = 2; act_sel_in[1] = 3; act_sel_in[2] = 1; act_sel_in[3] = 4; act_sel_in[4] = 3; act_sel_in[5] = 1; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 2; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 0; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=0; act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 1; act_sel_in[9] = 0; act_sel_in[10] = 0; act_sel_in[11] = 0; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 


#1.25 is_msb_in=1; column_idx_in=7; act[0] = -45; act[1] = 76; act[2] = -80; act[3] = 60; act[4] = 40; act[5] = 15; act[6] = 84; act[7] = -39; act[8] = -100; act[9] = -116; act[10] = -32; act[11] = 69; act[12] = -96; act[13] = -104; act[14] = 121; act[15] = -2; act[16] = 106; act[17] = 34; act[18] = 79; act[19] = 8; act[20] = 77; act[21] = -101; act[22] = -100; act[23] = -85; act[24] = -37; act[25] = -45; act[26] = 104; act[27] = -94; act[28] = -98; act[29] = 71; act[30] = -100; act[31] = -61; 
act_sel_in[0] = 0; act_sel_in[1] = 3; act_sel_in[2] = 4; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 4; act_sel_in[10] = 3; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 3; act_sel_in[14] = 3; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 is_msb_in=0; column_idx_in=6; act_sel_in[0] = 2; act_sel_in[1] = 3; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 2; act_sel_in[6] = 3; act_sel_in[7] = 0; act_sel_in[8] = 2; act_sel_in[9] = 0; act_sel_in[10] = 0; act_sel_in[11] = 3; act_sel_in[12] = 2; act_sel_in[13] = 3; act_sel_in[14] = 1; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=5; act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 2; act_sel_in[3] = 1; act_sel_in[4] = 3; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 2; act_sel_in[9] = 4; act_sel_in[10] = 0; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 1; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=4; act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 2; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 4; act_sel_in[6] = 3; act_sel_in[7] = 2; act_sel_in[8] = 3; act_sel_in[9] = 0; act_sel_in[10] = 3; act_sel_in[11] = 3; act_sel_in[12] = 3; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=3; act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 4; act_sel_in[9] = 0; act_sel_in[10] = 2; act_sel_in[11] = 0; act_sel_in[12] = 1; act_sel_in[13] = 3; act_sel_in[14] = 0; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=2; act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 4; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 4; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 2; act_sel_in[9] = 4; act_sel_in[10] = 3; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=1; act_sel_in[0] = 2; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 3; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 1; act_sel_in[7] = 3; act_sel_in[8] = 2; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 2; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 0; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=0; act_sel_in[0] = 1; act_sel_in[1] = 4; act_sel_in[2] = 4; act_sel_in[3] = 0; act_sel_in[4] = 0; act_sel_in[5] = 0; act_sel_in[6] = 4; act_sel_in[7] = 3; act_sel_in[8] = 1; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 0; act_sel_in[12] = 1; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 


#1.25 is_msb_in=1; column_idx_in=7; act[0] = 48; act[1] = -48; act[2] = 6; act[3] = -115; act[4] = 24; act[5] = 72; act[6] = 37; act[7] = 19; act[8] = 4; act[9] = 107; act[10] = 51; act[11] = 6; act[12] = -66; act[13] = -25; act[14] = -49; act[15] = 65; act[16] = -106; act[17] = -82; act[18] = 83; act[19] = -127; act[20] = 82; act[21] = 68; act[22] = 6; act[23] = -71; act[24] = -86; act[25] = -50; act[26] = 69; act[27] = 61; act[28] = 115; act[29] = -2; act[30] = 47; act[31] = -101; 
act_sel_in[0] = 4; act_sel_in[1] = 0; act_sel_in[2] = 4; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 0; act_sel_in[7] = 3; act_sel_in[8] = 3; act_sel_in[9] = 1; act_sel_in[10] = 3; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 0; act_sel_in[14] = 1; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 is_msb_in=0; column_idx_in=6; act_sel_in[0] = 1; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 2; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 1; act_sel_in[8] = 3; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 3; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=5; act_sel_in[0] = 0; act_sel_in[1] = 3; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 0; act_sel_in[8] = 4; act_sel_in[9] = 2; act_sel_in[10] = 1; act_sel_in[11] = 4; act_sel_in[12] = 1; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=4; act_sel_in[0] = 1; act_sel_in[1] = 0; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 4; act_sel_in[6] = 3; act_sel_in[7] = 2; act_sel_in[8] = 0; act_sel_in[9] = 2; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 3; act_sel_in[13] = 0; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=3; act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 1; act_sel_in[3] = 3; act_sel_in[4] = 2; act_sel_in[5] = 4; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 0; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 2; act_sel_in[14] = 1; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=2; act_sel_in[0] = 2; act_sel_in[1] = 3; act_sel_in[2] = 0; act_sel_in[3] = 0; act_sel_in[4] = 0; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 1; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 0; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=1; act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 3; act_sel_in[9] = 2; act_sel_in[10] = 1; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 3; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=0; act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 3; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 0; act_sel_in[7] = 1; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 0; act_sel_in[14] = 0; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 


#1.25 is_msb_in=1; column_idx_in=7; act[0] = -52; act[1] = -121; act[2] = 14; act[3] = 35; act[4] = -73; act[5] = 21; act[6] = 64; act[7] = -7; act[8] = -59; act[9] = 11; act[10] = -47; act[11] = -106; act[12] = 71; act[13] = 26; act[14] = 97; act[15] = 76; act[16] = -51; act[17] = -64; act[18] = 78; act[19] = -47; act[20] = 72; act[21] = -14; act[22] = -91; act[23] = -48; act[24] = -91; act[25] = -80; act[26] = -51; act[27] = -79; act[28] = -39; act[29] = 126; act[30] = -67; act[31] = -94; 
act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 4; act_sel_in[3] = 0; act_sel_in[4] = 0; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 is_msb_in=0; column_idx_in=6; act_sel_in[0] = 2; act_sel_in[1] = 4; act_sel_in[2] = 1; act_sel_in[3] = 3; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 1; act_sel_in[11] = 3; act_sel_in[12] = 2; act_sel_in[13] = 0; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=5; act_sel_in[0] = 1; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 4; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 0; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=4; act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 1; act_sel_in[3] = 4; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 4; act_sel_in[10] = 3; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 1; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=3; act_sel_in[0] = 2; act_sel_in[1] = 0; act_sel_in[2] = 3; act_sel_in[3] = 2; act_sel_in[4] = 3; act_sel_in[5] = 1; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 2; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=2; act_sel_in[0] = 4; act_sel_in[1] = 0; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 0; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 2; act_sel_in[10] = 0; act_sel_in[11] = 4; act_sel_in[12] = 4; act_sel_in[13] = 1; act_sel_in[14] = 0; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=1; act_sel_in[0] = 3; act_sel_in[1] = 2; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 2; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=0; act_sel_in[0] = 0; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 0; act_sel_in[5] = 1; act_sel_in[6] = 2; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 2; act_sel_in[10] = 3; act_sel_in[11] = 2; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 


#1.25 is_msb_in=1; column_idx_in=7; act[0] = 29; act[1] = -69; act[2] = 51; act[3] = 27; act[4] = 75; act[5] = -118; act[6] = 74; act[7] = -83; act[8] = 40; act[9] = 119; act[10] = -25; act[11] = 115; act[12] = 61; act[13] = 42; act[14] = -73; act[15] = 15; act[16] = -33; act[17] = 74; act[18] = 12; act[19] = -42; act[20] = -12; act[21] = 124; act[22] = 109; act[23] = -13; act[24] = 19; act[25] = 49; act[26] = -7; act[27] = -60; act[28] = -88; act[29] = 120; act[30] = 58; act[31] = 62; 
act_sel_in[0] = 2; act_sel_in[1] = 0; act_sel_in[2] = 4; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 0; act_sel_in[7] = 2; act_sel_in[8] = 3; act_sel_in[9] = 0; act_sel_in[10] = 3; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 2; act_sel_in[14] = 1; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 is_msb_in=0; column_idx_in=6; act_sel_in[0] = 0; act_sel_in[1] = 1; act_sel_in[2] = 2; act_sel_in[3] = 3; act_sel_in[4] = 2; act_sel_in[5] = 4; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 1; act_sel_in[9] = 3; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 3; act_sel_in[14] = 3; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=5; act_sel_in[0] = 2; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 0; act_sel_in[5] = 1; act_sel_in[6] = 3; act_sel_in[7] = 2; act_sel_in[8] = 1; act_sel_in[9] = 0; act_sel_in[10] = 4; act_sel_in[11] = 4; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 0; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=4; act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 0; act_sel_in[8] = 4; act_sel_in[9] = 3; act_sel_in[10] = 1; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=3; act_sel_in[0] = 4; act_sel_in[1] = 0; act_sel_in[2] = 2; act_sel_in[3] = 1; act_sel_in[4] = 0; act_sel_in[5] = 4; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 2; act_sel_in[14] = 0; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=2; act_sel_in[0] = 4; act_sel_in[1] = 0; act_sel_in[2] = 4; act_sel_in[3] = 2; act_sel_in[4] = 0; act_sel_in[5] = 0; act_sel_in[6] = 1; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 3; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 0; act_sel_in[14] = 4; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=1; act_sel_in[0] = 2; act_sel_in[1] = 0; act_sel_in[2] = 4; act_sel_in[3] = 2; act_sel_in[4] = 4; act_sel_in[5] = 4; act_sel_in[6] = 3; act_sel_in[7] = 0; act_sel_in[8] = 4; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=0; act_sel_in[0] = 0; act_sel_in[1] = 0; act_sel_in[2] = 0; act_sel_in[3] = 3; act_sel_in[4] = 0; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 4; act_sel_in[8] = 2; act_sel_in[9] = 0; act_sel_in[10] = 1; act_sel_in[11] = 3; act_sel_in[12] = 1; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 


#1.25 is_msb_in=1; column_idx_in=7; act[0] = -104; act[1] = -37; act[2] = -30; act[3] = -72; act[4] = -125; act[5] = -20; act[6] = 34; act[7] = -115; act[8] = 112; act[9] = -37; act[10] = -93; act[11] = 13; act[12] = -39; act[13] = 127; act[14] = 49; act[15] = 82; act[16] = -9; act[17] = -71; act[18] = -87; act[19] = -9; act[20] = 124; act[21] = 35; act[22] = -128; act[23] = -10; act[24] = 105; act[25] = 50; act[26] = -86; act[27] = -95; act[28] = 72; act[29] = -24; act[30] = 112; act[31] = 121; 
act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 3; act_sel_in[8] = 2; act_sel_in[9] = 4; act_sel_in[10] = 0; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 2; act_sel_in[14] = 0; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 is_msb_in=0; column_idx_in=6; act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 2; act_sel_in[3] = 3; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 2; act_sel_in[9] = 0; act_sel_in[10] = 4; act_sel_in[11] = 0; act_sel_in[12] = 3; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=5; act_sel_in[0] = 4; act_sel_in[1] = 1; act_sel_in[2] = 3; act_sel_in[3] = 2; act_sel_in[4] = 0; act_sel_in[5] = 1; act_sel_in[6] = 1; act_sel_in[7] = 3; act_sel_in[8] = 4; act_sel_in[9] = 3; act_sel_in[10] = 4; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=4; act_sel_in[0] = 3; act_sel_in[1] = 2; act_sel_in[2] = 1; act_sel_in[3] = 4; act_sel_in[4] = 2; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 3; act_sel_in[9] = 2; act_sel_in[10] = 1; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 2; act_sel_in[14] = 3; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=3; act_sel_in[0] = 3; act_sel_in[1] = 0; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 1; act_sel_in[6] = 0; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 2; act_sel_in[11] = 2; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=2; act_sel_in[0] = 3; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 1; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 3; act_sel_in[9] = 1; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 4; act_sel_in[13] = 3; act_sel_in[14] = 0; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=1; act_sel_in[0] = 3; act_sel_in[1] = 3; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 2; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 2; act_sel_in[9] = 0; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 3; act_sel_in[14] = 3; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=0; act_sel_in[0] = 0; act_sel_in[1] = 0; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 0; act_sel_in[5] = 4; act_sel_in[6] = 3; act_sel_in[7] = 2; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 


#1.25 is_msb_in=1; column_idx_in=7; act[0] = 7; act[1] = 56; act[2] = 43; act[3] = -68; act[4] = 31; act[5] = 3; act[6] = -102; act[7] = -43; act[8] = -68; act[9] = -106; act[10] = 21; act[11] = 82; act[12] = -33; act[13] = 98; act[14] = 18; act[15] = -82; act[16] = 112; act[17] = 49; act[18] = -27; act[19] = -93; act[20] = -12; act[21] = 116; act[22] = 97; act[23] = 109; act[24] = -112; act[25] = -119; act[26] = -72; act[27] = -107; act[28] = 98; act[29] = -43; act[30] = 100; act[31] = -95; 
act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 4; act_sel_in[9] = 0; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 is_msb_in=0; column_idx_in=6; act_sel_in[0] = 2; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 3; act_sel_in[4] = 0; act_sel_in[5] = 4; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 2; act_sel_in[9] = 3; act_sel_in[10] = 2; act_sel_in[11] = 0; act_sel_in[12] = 3; act_sel_in[13] = 4; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=5; act_sel_in[0] = 2; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 3; act_sel_in[11] = 3; act_sel_in[12] = 1; act_sel_in[13] = 2; act_sel_in[14] = 0; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=4; act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 2; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 1; act_sel_in[9] = 3; act_sel_in[10] = 0; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 3; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=3; act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 4; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 3; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 1; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=2; act_sel_in[0] = 4; act_sel_in[1] = 1; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 0; act_sel_in[7] = 1; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 4; act_sel_in[11] = 4; act_sel_in[12] = 1; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=1; act_sel_in[0] = 3; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 1; act_sel_in[7] = 1; act_sel_in[8] = 2; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 3; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 3; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=0; act_sel_in[0] = 4; act_sel_in[1] = 4; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 1; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 1; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 1; act_sel_in[12] = 2; act_sel_in[13] = 0; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 


#1.25 is_msb_in=1; column_idx_in=7; act[0] = 126; act[1] = 88; act[2] = 78; act[3] = 102; act[4] = -54; act[5] = -37; act[6] = -106; act[7] = 99; act[8] = 83; act[9] = -47; act[10] = -33; act[11] = -2; act[12] = 85; act[13] = 63; act[14] = 21; act[15] = 111; act[16] = -50; act[17] = 106; act[18] = 48; act[19] = 24; act[20] = 27; act[21] = 74; act[22] = 101; act[23] = 69; act[24] = -116; act[25] = 55; act[26] = 51; act[27] = -40; act[28] = 126; act[29] = 87; act[30] = -108; act[31] = -20; 
act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 0; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 0; act_sel_in[10] = 2; act_sel_in[11] = 0; act_sel_in[12] = 3; act_sel_in[13] = 3; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 is_msb_in=0; column_idx_in=6; act_sel_in[0] = 4; act_sel_in[1] = 3; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 2; act_sel_in[5] = 3; act_sel_in[6] = 2; act_sel_in[7] = 3; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=5; act_sel_in[0] = 2; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 3; act_sel_in[5] = 1; act_sel_in[6] = 2; act_sel_in[7] = 3; act_sel_in[8] = 1; act_sel_in[9] = 2; act_sel_in[10] = 1; act_sel_in[11] = 0; act_sel_in[12] = 4; act_sel_in[13] = 0; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=4; act_sel_in[0] = 4; act_sel_in[1] = 3; act_sel_in[2] = 3; act_sel_in[3] = 4; act_sel_in[4] = 0; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 1; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 2; act_sel_in[12] = 4; act_sel_in[13] = 0; act_sel_in[14] = 0; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=3; act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 4; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 3; act_sel_in[7] = 1; act_sel_in[8] = 3; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 2; act_sel_in[14] = 1; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=2; act_sel_in[0] = 4; act_sel_in[1] = 1; act_sel_in[2] = 0; act_sel_in[3] = 1; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 3; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 2; act_sel_in[14] = 1; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=1; act_sel_in[0] = 0; act_sel_in[1] = 0; act_sel_in[2] = 0; act_sel_in[3] = 3; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 4; act_sel_in[9] = 3; act_sel_in[10] = 3; act_sel_in[11] = 3; act_sel_in[12] = 1; act_sel_in[13] = 4; act_sel_in[14] = 2; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=0; act_sel_in[0] = 4; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 0; act_sel_in[4] = 0; act_sel_in[5] = 3; act_sel_in[6] = 1; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 0; act_sel_in[10] = 3; act_sel_in[11] = 3; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 3; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 


#1.25 is_msb_in=1; column_idx_in=7; act[0] = -12; act[1] = 33; act[2] = -96; act[3] = -9; act[4] = -28; act[5] = -47; act[6] = 65; act[7] = -27; act[8] = 55; act[9] = 14; act[10] = 56; act[11] = -122; act[12] = 114; act[13] = 14; act[14] = 53; act[15] = 71; act[16] = 96; act[17] = 70; act[18] = 14; act[19] = -81; act[20] = -22; act[21] = 48; act[22] = 41; act[23] = 18; act[24] = 92; act[25] = 113; act[26] = 46; act[27] = 69; act[28] = -40; act[29] = -46; act[30] = 75; act[31] = -9; 
act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 2; act_sel_in[3] = 3; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 2; act_sel_in[10] = 0; act_sel_in[11] = 0; act_sel_in[12] = 1; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 is_msb_in=0; column_idx_in=6; act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 3; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 3; act_sel_in[9] = 2; act_sel_in[10] = 2; act_sel_in[11] = 3; act_sel_in[12] = 1; act_sel_in[13] = 1; act_sel_in[14] = 1; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=5; act_sel_in[0] = 2; act_sel_in[1] = 2; act_sel_in[2] = 2; act_sel_in[3] = 1; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 4; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 0; act_sel_in[14] = 0; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=4; act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 2; act_sel_in[3] = 3; act_sel_in[4] = 0; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 4; act_sel_in[8] = 4; act_sel_in[9] = 2; act_sel_in[10] = 1; act_sel_in[11] = 3; act_sel_in[12] = 4; act_sel_in[13] = 3; act_sel_in[14] = 3; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=3; act_sel_in[0] = 1; act_sel_in[1] = 1; act_sel_in[2] = 4; act_sel_in[3] = 3; act_sel_in[4] = 2; act_sel_in[5] = 1; act_sel_in[6] = 2; act_sel_in[7] = 2; act_sel_in[8] = 1; act_sel_in[9] = 1; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 2; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=2; act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 4; act_sel_in[6] = 1; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 3; act_sel_in[12] = 3; act_sel_in[13] = 3; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=1; act_sel_in[0] = 2; act_sel_in[1] = 3; act_sel_in[2] = 4; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 1; act_sel_in[7] = 1; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 3; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=0; act_sel_in[0] = 0; act_sel_in[1] = 3; act_sel_in[2] = 3; act_sel_in[3] = 2; act_sel_in[4] = 2; act_sel_in[5] = 3; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 3; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 


#1.25 is_msb_in=1; column_idx_in=7; act[0] = -18; act[1] = -81; act[2] = 35; act[3] = -93; act[4] = -60; act[5] = 58; act[6] = 45; act[7] = 7; act[8] = -22; act[9] = -20; act[10] = -36; act[11] = 6; act[12] = 19; act[13] = 117; act[14] = -81; act[15] = -100; act[16] = -40; act[17] = 43; act[18] = 89; act[19] = 94; act[20] = 16; act[21] = -106; act[22] = 122; act[23] = 41; act[24] = -111; act[25] = -119; act[26] = -3; act[27] = 83; act[28] = 56; act[29] = 68; act[30] = 34; act[31] = 80; 
act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 4; act_sel_in[11] = 0; act_sel_in[12] = 3; act_sel_in[13] = 1; act_sel_in[14] = 3; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 is_msb_in=0; column_idx_in=6; act_sel_in[0] = 1; act_sel_in[1] = 0; act_sel_in[2] = 0; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 3; act_sel_in[8] = 2; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 4; act_sel_in[12] = 4; act_sel_in[13] = 3; act_sel_in[14] = 0; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=5; act_sel_in[0] = 0; act_sel_in[1] = 3; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 3; act_sel_in[5] = 4; act_sel_in[6] = 0; act_sel_in[7] = 2; act_sel_in[8] = 1; act_sel_in[9] = 2; act_sel_in[10] = 2; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 4; act_sel_in[14] = 1; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=4; act_sel_in[0] = 2; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 1; act_sel_in[6] = 3; act_sel_in[7] = 2; act_sel_in[8] = 4; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 4; act_sel_in[12] = 4; act_sel_in[13] = 3; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=3; act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 2; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 2; act_sel_in[11] = 2; act_sel_in[12] = 4; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=2; act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 0; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 4; act_sel_in[9] = 3; act_sel_in[10] = 4; act_sel_in[11] = 3; act_sel_in[12] = 3; act_sel_in[13] = 1; act_sel_in[14] = 3; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=1; act_sel_in[0] = 4; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 0; act_sel_in[6] = 4; act_sel_in[7] = 4; act_sel_in[8] = 4; act_sel_in[9] = 0; act_sel_in[10] = 0; act_sel_in[11] = 2; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 1; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=0; act_sel_in[0] = 2; act_sel_in[1] = 3; act_sel_in[2] = 3; act_sel_in[3] = 2; act_sel_in[4] = 0; act_sel_in[5] = 3; act_sel_in[6] = 4; act_sel_in[7] = 4; act_sel_in[8] = 2; act_sel_in[9] = 3; act_sel_in[10] = 0; act_sel_in[11] = 4; act_sel_in[12] = 4; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 


#1.25 is_msb_in=1; column_idx_in=7; act[0] = -42; act[1] = 109; act[2] = 88; act[3] = -127; act[4] = -83; act[5] = 46; act[6] = 93; act[7] = -81; act[8] = -53; act[9] = 0; act[10] = 120; act[11] = 80; act[12] = 27; act[13] = 18; act[14] = 59; act[15] = -78; act[16] = -43; act[17] = -48; act[18] = -67; act[19] = -70; act[20] = 45; act[21] = -98; act[22] = -110; act[23] = 63; act[24] = -12; act[25] = -105; act[26] = -22; act[27] = 99; act[28] = -52; act[29] = 55; act[30] = 84; act[31] = 72; 
act_sel_in[0] = 3; act_sel_in[1] = 0; act_sel_in[2] = 4; act_sel_in[3] = 4; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 0; act_sel_in[7] = 1; act_sel_in[8] = 2; act_sel_in[9] = 0; act_sel_in[10] = 2; act_sel_in[11] = 0; act_sel_in[12] = 4; act_sel_in[13] = 4; act_sel_in[14] = 1; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 is_msb_in=0; column_idx_in=6; act_sel_in[0] = 2; act_sel_in[1] = 4; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 3; act_sel_in[8] = 3; act_sel_in[9] = 4; act_sel_in[10] = 3; act_sel_in[11] = 0; act_sel_in[12] = 1; act_sel_in[13] = 1; act_sel_in[14] = 0; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=5; act_sel_in[0] = 3; act_sel_in[1] = 3; act_sel_in[2] = 3; act_sel_in[3] = 4; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 3; act_sel_in[9] = 1; act_sel_in[10] = 4; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=4; act_sel_in[0] = 0; act_sel_in[1] = 3; act_sel_in[2] = 4; act_sel_in[3] = 1; act_sel_in[4] = 3; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 2; act_sel_in[8] = 4; act_sel_in[9] = 0; act_sel_in[10] = 1; act_sel_in[11] = 4; act_sel_in[12] = 4; act_sel_in[13] = 0; act_sel_in[14] = 3; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=3; act_sel_in[0] = 0; act_sel_in[1] = 1; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 0; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 2; act_sel_in[8] = 2; act_sel_in[9] = 4; act_sel_in[10] = 3; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 1; act_sel_in[14] = 0; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=2; act_sel_in[0] = 4; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 0; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 2; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 2; act_sel_in[14] = 3; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=1; act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 4; act_sel_in[11] = 0; act_sel_in[12] = 4; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=0; act_sel_in[0] = 4; act_sel_in[1] = 4; act_sel_in[2] = 0; act_sel_in[3] = 1; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 


#1.25 is_msb_in=1; column_idx_in=7; act[0] = 88; act[1] = 52; act[2] = 104; act[3] = 89; act[4] = -65; act[5] = 55; act[6] = -113; act[7] = -21; act[8] = -43; act[9] = 70; act[10] = 5; act[11] = -61; act[12] = 79; act[13] = -63; act[14] = -99; act[15] = 100; act[16] = 117; act[17] = -125; act[18] = -30; act[19] = -122; act[20] = 99; act[21] = 109; act[22] = 64; act[23] = -78; act[24] = -109; act[25] = -108; act[26] = 14; act[27] = -61; act[28] = -36; act[29] = 102; act[30] = 101; act[31] = -22; 
act_sel_in[0] = 3; act_sel_in[1] = 2; act_sel_in[2] = 4; act_sel_in[3] = 1; act_sel_in[4] = 3; act_sel_in[5] = 4; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 2; act_sel_in[13] = 0; act_sel_in[14] = 3; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 is_msb_in=0; column_idx_in=6; act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 4; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 2; act_sel_in[7] = 3; act_sel_in[8] = 3; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 4; act_sel_in[12] = 1; act_sel_in[13] = 2; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=5; act_sel_in[0] = 1; act_sel_in[1] = 0; act_sel_in[2] = 0; act_sel_in[3] = 2; act_sel_in[4] = 0; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 2; act_sel_in[9] = 4; act_sel_in[10] = 4; act_sel_in[11] = 4; act_sel_in[12] = 4; act_sel_in[13] = 3; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=4; act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 0; act_sel_in[10] = 3; act_sel_in[11] = 3; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=3; act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 4; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 4; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 4; act_sel_in[12] = 1; act_sel_in[13] = 0; act_sel_in[14] = 1; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=2; act_sel_in[0] = 4; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 3; act_sel_in[5] = 4; act_sel_in[6] = 1; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 0; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 3; act_sel_in[13] = 3; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=1; act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 2; act_sel_in[5] = 4; act_sel_in[6] = 4; act_sel_in[7] = 0; act_sel_in[8] = 3; act_sel_in[9] = 1; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 1; act_sel_in[14] = 1; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=0; act_sel_in[0] = 3; act_sel_in[1] = 1; act_sel_in[2] = 0; act_sel_in[3] = 1; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 3; act_sel_in[8] = 2; act_sel_in[9] = 3; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 2; act_sel_in[13] = 0; act_sel_in[14] = 3; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 


#1.25 is_msb_in=1; column_idx_in=7; act[0] = -4; act[1] = 95; act[2] = -103; act[3] = -115; act[4] = 24; act[5] = 70; act[6] = -75; act[7] = 73; act[8] = 108; act[9] = -87; act[10] = -95; act[11] = -104; act[12] = 108; act[13] = 80; act[14] = -119; act[15] = -1; act[16] = -102; act[17] = -12; act[18] = -54; act[19] = -20; act[20] = 10; act[21] = -38; act[22] = 30; act[23] = 59; act[24] = 51; act[25] = -27; act[26] = 44; act[27] = 92; act[28] = -120; act[29] = -104; act[30] = 31; act[31] = -127; 
act_sel_in[0] = 0; act_sel_in[1] = 1; act_sel_in[2] = 0; act_sel_in[3] = 3; act_sel_in[4] = 3; act_sel_in[5] = 4; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 1; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 1; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 3; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 is_msb_in=0; column_idx_in=6; act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 0; act_sel_in[10] = 0; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 0; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=5; act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 1; act_sel_in[7] = 1; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 0; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=4; act_sel_in[0] = 3; act_sel_in[1] = 0; act_sel_in[2] = 2; act_sel_in[3] = 3; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 3; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 1; act_sel_in[10] = 4; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=3; act_sel_in[0] = 4; act_sel_in[1] = 1; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 1; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 3; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 0; act_sel_in[14] = 1; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=2; act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 0; act_sel_in[5] = 0; act_sel_in[6] = 0; act_sel_in[7] = 3; act_sel_in[8] = 2; act_sel_in[9] = 1; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 3; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=1; act_sel_in[0] = 2; act_sel_in[1] = 2; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 0; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 3; act_sel_in[12] = 4; act_sel_in[13] = 0; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=0; act_sel_in[0] = 0; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 1; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 1; act_sel_in[11] = 3; act_sel_in[12] = 4; act_sel_in[13] = 0; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 


#1.25 is_msb_in=1; column_idx_in=7; act[0] = -46; act[1] = 103; act[2] = -78; act[3] = 8; act[4] = -68; act[5] = 37; act[6] = 7; act[7] = -17; act[8] = -40; act[9] = 106; act[10] = 43; act[11] = 7; act[12] = -89; act[13] = -73; act[14] = -67; act[15] = 10; act[16] = 76; act[17] = 4; act[18] = 100; act[19] = -31; act[20] = -86; act[21] = 77; act[22] = -109; act[23] = 57; act[24] = 108; act[25] = 21; act[26] = -42; act[27] = -22; act[28] = -94; act[29] = -104; act[30] = -44; act[31] = 30; 
act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 1; act_sel_in[3] = 3; act_sel_in[4] = 4; act_sel_in[5] = 4; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 3; act_sel_in[14] = 3; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 is_msb_in=0; column_idx_in=6; act_sel_in[0] = 0; act_sel_in[1] = 1; act_sel_in[2] = 4; act_sel_in[3] = 4; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 1; act_sel_in[9] = 0; act_sel_in[10] = 1; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 3; act_sel_in[14] = 4; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=5; act_sel_in[0] = 2; act_sel_in[1] = 0; act_sel_in[2] = 2; act_sel_in[3] = 3; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 0; act_sel_in[9] = 2; act_sel_in[10] = 0; act_sel_in[11] = 3; act_sel_in[12] = 4; act_sel_in[13] = 3; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=4; act_sel_in[0] = 1; act_sel_in[1] = 0; act_sel_in[2] = 4; act_sel_in[3] = 2; act_sel_in[4] = 3; act_sel_in[5] = 1; act_sel_in[6] = 1; act_sel_in[7] = 4; act_sel_in[8] = 1; act_sel_in[9] = 0; act_sel_in[10] = 0; act_sel_in[11] = 4; act_sel_in[12] = 1; act_sel_in[13] = 4; act_sel_in[14] = 3; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=3; act_sel_in[0] = 4; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 3; act_sel_in[6] = 4; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 4; act_sel_in[10] = 4; act_sel_in[11] = 3; act_sel_in[12] = 3; act_sel_in[13] = 4; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=2; act_sel_in[0] = 3; act_sel_in[1] = 3; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 3; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 3; act_sel_in[13] = 0; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=1; act_sel_in[0] = 2; act_sel_in[1] = 2; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 1; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 2; act_sel_in[8] = 2; act_sel_in[9] = 4; act_sel_in[10] = 4; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 2; act_sel_in[14] = 1; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=0; act_sel_in[0] = 1; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 4; act_sel_in[4] = 2; act_sel_in[5] = 1; act_sel_in[6] = 2; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 0; act_sel_in[12] = 3; act_sel_in[13] = 1; act_sel_in[14] = 3; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 


#1.25 is_msb_in=1; column_idx_in=7; act[0] = -18; act[1] = 94; act[2] = 14; act[3] = -54; act[4] = 68; act[5] = -100; act[6] = -53; act[7] = -61; act[8] = -97; act[9] = 63; act[10] = -11; act[11] = -63; act[12] = 81; act[13] = 3; act[14] = 94; act[15] = -72; act[16] = 23; act[17] = 40; act[18] = 86; act[19] = 88; act[20] = -88; act[21] = -111; act[22] = -64; act[23] = 111; act[24] = 29; act[25] = -24; act[26] = -7; act[27] = -106; act[28] = -5; act[29] = 109; act[30] = -116; act[31] = 53; 
act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 2; act_sel_in[7] = 2; act_sel_in[8] = 4; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 3; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 1; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 is_msb_in=0; column_idx_in=6; act_sel_in[0] = 3; act_sel_in[1] = 0; act_sel_in[2] = 1; act_sel_in[3] = 3; act_sel_in[4] = 4; act_sel_in[5] = 4; act_sel_in[6] = 4; act_sel_in[7] = 3; act_sel_in[8] = 2; act_sel_in[9] = 0; act_sel_in[10] = 3; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=5; act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 1; act_sel_in[4] = 1; act_sel_in[5] = 4; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 2; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 4; act_sel_in[12] = 1; act_sel_in[13] = 0; act_sel_in[14] = 0; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=4; act_sel_in[0] = 4; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 0; act_sel_in[5] = 0; act_sel_in[6] = 1; act_sel_in[7] = 4; act_sel_in[8] = 4; act_sel_in[9] = 2; act_sel_in[10] = 3; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=3; act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 0; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 4; act_sel_in[6] = 0; act_sel_in[7] = 1; act_sel_in[8] = 1; act_sel_in[9] = 0; act_sel_in[10] = 1; act_sel_in[11] = 4; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=2; act_sel_in[0] = 4; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 2; act_sel_in[5] = 2; act_sel_in[6] = 0; act_sel_in[7] = 1; act_sel_in[8] = 2; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 3; act_sel_in[14] = 1; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=1; act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 2; act_sel_in[3] = 2; act_sel_in[4] = 3; act_sel_in[5] = 4; act_sel_in[6] = 3; act_sel_in[7] = 1; act_sel_in[8] = 0; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 3; act_sel_in[12] = 3; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=0; act_sel_in[0] = 3; act_sel_in[1] = 3; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 2; act_sel_in[10] = 2; act_sel_in[11] = 2; act_sel_in[12] = 3; act_sel_in[13] = 2; act_sel_in[14] = 3; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 


#1.25 is_msb_in=1; column_idx_in=7; act[0] = 113; act[1] = -11; act[2] = -38; act[3] = 12; act[4] = -126; act[5] = -19; act[6] = -46; act[7] = 109; act[8] = -119; act[9] = -24; act[10] = -2; act[11] = 63; act[12] = -27; act[13] = 66; act[14] = 127; act[15] = -43; act[16] = -78; act[17] = -43; act[18] = 96; act[19] = -117; act[20] = 18; act[21] = 116; act[22] = -41; act[23] = -83; act[24] = -94; act[25] = -46; act[26] = -94; act[27] = 93; act[28] = -41; act[29] = 89; act[30] = 73; act[31] = 104; 
act_sel_in[0] = 0; act_sel_in[1] = 3; act_sel_in[2] = 3; act_sel_in[3] = 2; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 2; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 1; act_sel_in[11] = 4; act_sel_in[12] = 3; act_sel_in[13] = 4; act_sel_in[14] = 3; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 is_msb_in=0; column_idx_in=6; act_sel_in[0] = 3; act_sel_in[1] = 0; act_sel_in[2] = 3; act_sel_in[3] = 2; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 4; act_sel_in[9] = 3; act_sel_in[10] = 2; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 4; act_sel_in[14] = 3; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=5; act_sel_in[0] = 1; act_sel_in[1] = 1; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 4; act_sel_in[5] = 4; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 3; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 4; act_sel_in[14] = 2; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=4; act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 0; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 4; act_sel_in[9] = 0; act_sel_in[10] = 4; act_sel_in[11] = 0; act_sel_in[12] = 3; act_sel_in[13] = 0; act_sel_in[14] = 1; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=3; act_sel_in[0] = 4; act_sel_in[1] = 4; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 2; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 3; act_sel_in[11] = 1; act_sel_in[12] = 0; act_sel_in[13] = 4; act_sel_in[14] = 1; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=2; act_sel_in[0] = 2; act_sel_in[1] = 2; act_sel_in[2] = 1; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 4; act_sel_in[9] = 4; act_sel_in[10] = 3; act_sel_in[11] = 2; act_sel_in[12] = 0; act_sel_in[13] = 4; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=1; act_sel_in[0] = 2; act_sel_in[1] = 2; act_sel_in[2] = 4; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 2; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 3; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 2; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=0; act_sel_in[0] = 4; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 3; act_sel_in[4] = 0; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 1; act_sel_in[10] = 1; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 


#1.25 is_msb_in=1; column_idx_in=7; act[0] = 114; act[1] = -86; act[2] = 29; act[3] = -85; act[4] = -38; act[5] = 75; act[6] = -55; act[7] = 99; act[8] = 46; act[9] = -82; act[10] = 91; act[11] = -5; act[12] = -51; act[13] = 2; act[14] = 29; act[15] = 120; act[16] = 21; act[17] = -121; act[18] = 43; act[19] = -98; act[20] = -34; act[21] = 112; act[22] = 39; act[23] = -85; act[24] = 101; act[25] = 116; act[26] = 121; act[27] = 68; act[28] = -97; act[29] = 125; act[30] = -105; act[31] = 120; 
act_sel_in[0] = 0; act_sel_in[1] = 3; act_sel_in[2] = 0; act_sel_in[3] = 2; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 4; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 is_msb_in=0; column_idx_in=6; act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 0; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 3; act_sel_in[9] = 2; act_sel_in[10] = 3; act_sel_in[11] = 3; act_sel_in[12] = 4; act_sel_in[13] = 1; act_sel_in[14] = 3; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=5; act_sel_in[0] = 2; act_sel_in[1] = 3; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 0; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 4; act_sel_in[9] = 4; act_sel_in[10] = 3; act_sel_in[11] = 3; act_sel_in[12] = 1; act_sel_in[13] = 4; act_sel_in[14] = 1; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=4; act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 1; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 4; act_sel_in[6] = 2; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 1; act_sel_in[10] = 3; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 3; act_sel_in[14] = 3; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=3; act_sel_in[0] = 2; act_sel_in[1] = 0; act_sel_in[2] = 4; act_sel_in[3] = 3; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 0; act_sel_in[8] = 3; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 4; act_sel_in[12] = 3; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=2; act_sel_in[0] = 2; act_sel_in[1] = 3; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 2; act_sel_in[5] = 4; act_sel_in[6] = 3; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 0; act_sel_in[10] = 4; act_sel_in[11] = 2; act_sel_in[12] = 0; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=1; act_sel_in[0] = 3; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 2; act_sel_in[4] = 3; act_sel_in[5] = 1; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 2; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=0; act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 0; act_sel_in[5] = 1; act_sel_in[6] = 1; act_sel_in[7] = 3; act_sel_in[8] = 3; act_sel_in[9] = 2; act_sel_in[10] = 1; act_sel_in[11] = 3; act_sel_in[12] = 1; act_sel_in[13] = 4; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 


#1.25 is_msb_in=1; column_idx_in=7; act[0] = 70; act[1] = 16; act[2] = -30; act[3] = 13; act[4] = -42; act[5] = 94; act[6] = 7; act[7] = 91; act[8] = -71; act[9] = -46; act[10] = -82; act[11] = 68; act[12] = 120; act[13] = 21; act[14] = 119; act[15] = 1; act[16] = 93; act[17] = -77; act[18] = -33; act[19] = -50; act[20] = -30; act[21] = -10; act[22] = 83; act[23] = -87; act[24] = 101; act[25] = -80; act[26] = -124; act[27] = 95; act[28] = -72; act[29] = 110; act[30] = -92; act[31] = 42; 
act_sel_in[0] = 1; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 2; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 1; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 0; act_sel_in[14] = 1; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 is_msb_in=0; column_idx_in=6; act_sel_in[0] = 1; act_sel_in[1] = 4; act_sel_in[2] = 0; act_sel_in[3] = 0; act_sel_in[4] = 0; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 0; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 1; act_sel_in[11] = 0; act_sel_in[12] = 3; act_sel_in[13] = 3; act_sel_in[14] = 1; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=5; act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 3; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=4; act_sel_in[0] = 1; act_sel_in[1] = 4; act_sel_in[2] = 4; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 4; act_sel_in[11] = 4; act_sel_in[12] = 4; act_sel_in[13] = 4; act_sel_in[14] = 1; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=3; act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 0; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 4; act_sel_in[7] = 0; act_sel_in[8] = 2; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 0; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=2; act_sel_in[0] = 3; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 4; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 4; act_sel_in[10] = 3; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 1; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=1; act_sel_in[0] = 2; act_sel_in[1] = 2; act_sel_in[2] = 4; act_sel_in[3] = 0; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 2; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 4; act_sel_in[14] = 4; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=0; act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 4; act_sel_in[6] = 2; act_sel_in[7] = 3; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 2; act_sel_in[12] = 3; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 


#1.25 is_msb_in=1; column_idx_in=7; act[0] = 0; act[1] = 73; act[2] = 55; act[3] = -83; act[4] = -103; act[5] = -52; act[6] = 54; act[7] = -85; act[8] = -49; act[9] = 58; act[10] = -117; act[11] = 55; act[12] = -53; act[13] = 73; act[14] = 29; act[15] = 109; act[16] = 83; act[17] = -24; act[18] = 103; act[19] = -107; act[20] = -59; act[21] = 54; act[22] = -7; act[23] = -97; act[24] = -98; act[25] = 119; act[26] = 6; act[27] = 63; act[28] = 40; act[29] = 73; act[30] = 59; act[31] = -80; 
act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 3; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 3; act_sel_in[9] = 0; act_sel_in[10] = 0; act_sel_in[11] = 0; act_sel_in[12] = 1; act_sel_in[13] = 2; act_sel_in[14] = 0; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 is_msb_in=0; column_idx_in=6; act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 0; act_sel_in[7] = 2; act_sel_in[8] = 4; act_sel_in[9] = 3; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 0; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=5; act_sel_in[0] = 1; act_sel_in[1] = 0; act_sel_in[2] = 4; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 4; act_sel_in[6] = 0; act_sel_in[7] = 0; act_sel_in[8] = 3; act_sel_in[9] = 2; act_sel_in[10] = 2; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 0; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=4; act_sel_in[0] = 3; act_sel_in[1] = 2; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 2; act_sel_in[6] = 0; act_sel_in[7] = 3; act_sel_in[8] = 1; act_sel_in[9] = 1; act_sel_in[10] = 4; act_sel_in[11] = 3; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 0; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=3; act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 4; act_sel_in[3] = 0; act_sel_in[4] = 2; act_sel_in[5] = 4; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 1; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=2; act_sel_in[0] = 2; act_sel_in[1] = 3; act_sel_in[2] = 3; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 0; act_sel_in[14] = 1; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=1; act_sel_in[0] = 3; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 0; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 1; act_sel_in[12] = 0; act_sel_in[13] = 2; act_sel_in[14] = 1; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=0; act_sel_in[0] = 0; act_sel_in[1] = 0; act_sel_in[2] = 3; act_sel_in[3] = 2; act_sel_in[4] = 0; act_sel_in[5] = 3; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 3; act_sel_in[10] = 0; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 4; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 


#1.25 is_msb_in=1; column_idx_in=7; act[0] = 93; act[1] = 112; act[2] = -14; act[3] = 44; act[4] = 57; act[5] = 32; act[6] = 108; act[7] = 63; act[8] = 77; act[9] = -25; act[10] = 50; act[11] = -75; act[12] = 91; act[13] = 69; act[14] = 70; act[15] = -22; act[16] = -38; act[17] = -13; act[18] = 1; act[19] = -123; act[20] = 48; act[21] = 4; act[22] = 32; act[23] = -114; act[24] = -78; act[25] = -18; act[26] = 102; act[27] = -98; act[28] = -63; act[29] = 54; act[30] = 26; act[31] = -82; 
act_sel_in[0] = 4; act_sel_in[1] = 0; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 2; act_sel_in[5] = 3; act_sel_in[6] = 1; act_sel_in[7] = 1; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 0; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 is_msb_in=0; column_idx_in=6; act_sel_in[0] = 1; act_sel_in[1] = 0; act_sel_in[2] = 0; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=5; act_sel_in[0] = 4; act_sel_in[1] = 3; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 2; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 4; act_sel_in[12] = 1; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=4; act_sel_in[0] = 4; act_sel_in[1] = 0; act_sel_in[2] = 4; act_sel_in[3] = 3; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 2; act_sel_in[8] = 1; act_sel_in[9] = 0; act_sel_in[10] = 4; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=3; act_sel_in[0] = 3; act_sel_in[1] = 0; act_sel_in[2] = 2; act_sel_in[3] = 0; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 3; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 0; act_sel_in[14] = 4; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=2; act_sel_in[0] = 4; act_sel_in[1] = 0; act_sel_in[2] = 2; act_sel_in[3] = 0; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 4; act_sel_in[9] = 2; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 4; act_sel_in[14] = 1; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=1; act_sel_in[0] = 3; act_sel_in[1] = 3; act_sel_in[2] = 4; act_sel_in[3] = 1; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 2; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 4; act_sel_in[12] = 1; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=0; act_sel_in[0] = 3; act_sel_in[1] = 2; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 0; act_sel_in[7] = 0; act_sel_in[8] = 2; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 0; act_sel_in[14] = 3; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 


#1.25 is_msb_in=1; column_idx_in=7; act[0] = 104; act[1] = -105; act[2] = -5; act[3] = 25; act[4] = -42; act[5] = 109; act[6] = -36; act[7] = 0; act[8] = 61; act[9] = 117; act[10] = -17; act[11] = -94; act[12] = 44; act[13] = -33; act[14] = -108; act[15] = -89; act[16] = -93; act[17] = 85; act[18] = -108; act[19] = 124; act[20] = -6; act[21] = -90; act[22] = -1; act[23] = -65; act[24] = 119; act[25] = 62; act[26] = 42; act[27] = -94; act[28] = 51; act[29] = -43; act[30] = -109; act[31] = -45; 
act_sel_in[0] = 1; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 2; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 1; act_sel_in[7] = 3; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 4; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 0; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 is_msb_in=0; column_idx_in=6; act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 4; act_sel_in[3] = 1; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 4; act_sel_in[8] = 4; act_sel_in[9] = 2; act_sel_in[10] = 2; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=5; act_sel_in[0] = 2; act_sel_in[1] = 3; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 2; act_sel_in[6] = 0; act_sel_in[7] = 3; act_sel_in[8] = 1; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=4; act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 0; act_sel_in[5] = 0; act_sel_in[6] = 0; act_sel_in[7] = 0; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 1; act_sel_in[11] = 0; act_sel_in[12] = 3; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=3; act_sel_in[0] = 0; act_sel_in[1] = 3; act_sel_in[2] = 4; act_sel_in[3] = 0; act_sel_in[4] = 2; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 3; act_sel_in[8] = 1; act_sel_in[9] = 3; act_sel_in[10] = 3; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=2; act_sel_in[0] = 2; act_sel_in[1] = 4; act_sel_in[2] = 4; act_sel_in[3] = 2; act_sel_in[4] = 4; act_sel_in[5] = 4; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 1; act_sel_in[9] = 3; act_sel_in[10] = 0; act_sel_in[11] = 0; act_sel_in[12] = 4; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 1; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 1; 
#1.25 column_idx_in=1; act_sel_in[0] = 2; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 3; act_sel_in[5] = 0; act_sel_in[6] = 0; act_sel_in[7] = 4; act_sel_in[8] = 1; act_sel_in[9] = 0; act_sel_in[10] = 0; act_sel_in[11] = 0; act_sel_in[12] = 3; act_sel_in[13] = 1; act_sel_in[14] = 3; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero_in[0] = 0; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 0; is_skip_zero_in[3] = 0; 
#1.25 column_idx_in=0; act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 3; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 4; act_sel_in[6] = 0; act_sel_in[7] = 1; act_sel_in[8] = 4; act_sel_in[9] = 0; act_sel_in[10] = 4; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 0; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero_in[0] = 1; is_skip_zero_in[1] = 0; is_skip_zero_in[2] = 1; is_skip_zero_in[3] = 1; 






    #15 $stop;
  end

  always #1.25 clk = ~clk;

endmodule

`endif