`ifndef __vert_32_tb_V__
`define __vert_32_tb_V__

`include "mac_unit_Vert_32_no_mul.v"

module vert_32_tb;
    
    parameter DATA_WIDTH    = 8;
    parameter VEC_LENGTH    = 32;
    parameter MUX_SEL_WIDTH = 3;
    parameter SUM_ACT_WIDTH = $clog2(VEC_LENGTH) + DATA_WIDTH - 2;
    parameter ACC_WIDTH     = DATA_WIDTH + 16;
    parameter RESULT_WIDTH  = 2*DATA_WIDTH;

    logic                               clk;
	logic                               reset;
	logic                               en_acc;
	logic                               load_accum;

	logic signed   [DATA_WIDTH-1:0]     act_in   [VEC_LENGTH-1:0];   // input activation (signed)
	logic          [MUX_SEL_WIDTH-1:0]  act_sel_in  [VEC_LENGTH/2-1:0]; // input activation MUX select signal
	logic                               act_val_in  [VEC_LENGTH/2-1:0]; // whether activation is valid
	logic signed   [SUM_ACT_WIDTH-1:0]  sum_act  [VEC_LENGTH/8-1:0]; // sum of a group of activations (signed)

	logic          [2:0]                column_idx;    // current column index for shifting 
	logic                               is_msb;        // specify if the current column is MSB
	logic                               is_skip_zero [VEC_LENGTH/8-1:0];  // specify if skip bit 0
	
	logic signed   [ACC_WIDTH-1:0]      accum_prev;
    logic signed   [RESULT_WIDTH-1:0]   result;

    mac_unit_Vert_32_no_mul_clk #(DATA_WIDTH, VEC_LENGTH, MUX_SEL_WIDTH, SUM_ACT_WIDTH, ACC_WIDTH) s (.*);

  initial
    $monitor ("out=%b", result);

  initial begin
    #0 clk = 0; reset = 1;  en_acc = 0;
    #1.2 reset = 0; en_acc = 1; load_accum = 0; accum_prev = 0;

    #1 is_msb=1; column_idx=7; act_in[0] = -50; act_in[1] = -79; act_in[2] = 6; act_in[3] = -2; act_in[4] = 100; act_in[5] = 74; act_in[6] = -9; act_in[7] = -88; act_in[8] = 38; act_in[9] = -44; act_in[10] = -90; act_in[11] = -77; act_in[12] = 4; act_in[13] = 10; act_in[14] = 83; act_in[15] = -100; act_in[16] = -83; act_in[17] = 122; act_in[18] = 25; act_in[19] = 93; act_in[20] = 97; act_in[21] = -79; act_in[22] = 30; act_in[23] = 53; act_in[24] = -61; act_in[25] = 1; act_in[26] = 76; act_in[27] = -127; act_in[28] = -49; act_in[29] = 102; act_in[30] = -18; act_in[31] = -57; 
    act_sel_in[0] = 3; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 3; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 1; act_sel_in[9] = 4; act_sel_in[10] = 3; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 2; act_sel_in[1] = 2; act_sel_in[2] = 2; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 4; act_sel_in[6] = 4; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 4; act_sel_in[14] = 4; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=5; act_sel_in[0] = 4; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 4; act_sel_in[9] = 0; act_sel_in[10] = 4; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=4; act_sel_in[0] = 1; act_sel_in[1] = 0; act_sel_in[2] = 2; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 0; act_sel_in[7] = 2; act_sel_in[8] = 1; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 2; act_sel_in[12] = 3; act_sel_in[13] = 4; act_sel_in[14] = 3; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 0; act_sel_in[1] = 1; act_sel_in[2] = 2; act_sel_in[3] = 0; act_sel_in[4] = 4; act_sel_in[5] = 4; act_sel_in[6] = 2; act_sel_in[7] = 2; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 3; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 1; act_sel_in[14] = 1; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=2; act_sel_in[0] = 0; act_sel_in[1] = 3; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 3; act_sel_in[6] = 0; act_sel_in[7] = 1; act_sel_in[8] = 4; act_sel_in[9] = 3; act_sel_in[10] = 1; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 2; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=1; act_sel_in[0] = 3; act_sel_in[1] = 3; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 2; act_sel_in[8] = 1; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=0; act_sel_in[0] = 0; act_sel_in[1] = 1; act_sel_in[2] = 0; act_sel_in[3] = 3; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 0; act_sel_in[7] = 1; act_sel_in[8] = 1; act_sel_in[9] = 2; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 0; act_sel_in[13] = 0; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 


    #1 is_msb=1; column_idx=7; act_in[0] = -49; act_in[1] = 49; act_in[2] = -84; act_in[3] = -93; act_in[4] = -126; act_in[5] = -72; act_in[6] = 56; act_in[7] = -28; act_in[8] = 10; act_in[9] = 15; act_in[10] = 28; act_in[11] = 90; act_in[12] = -91; act_in[13] = 125; act_in[14] = 0; act_in[15] = 5; act_in[16] = 6; act_in[17] = -20; act_in[18] = -26; act_in[19] = -17; act_in[20] = -98; act_in[21] = -115; act_in[22] = -117; act_in[23] = 0; act_in[24] = 16; act_in[25] = 125; act_in[26] = -23; act_in[27] = 54; act_in[28] = -58; act_in[29] = -60; act_in[30] = -8; act_in[31] = 61; 
    act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 4; act_sel_in[3] = 2; act_sel_in[4] = 4; act_sel_in[5] = 4; act_sel_in[6] = 1; act_sel_in[7] = 1; act_sel_in[8] = 3; act_sel_in[9] = 0; act_sel_in[10] = 2; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 1; act_sel_in[14] = 0; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 2; act_sel_in[1] = 4; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 2; act_sel_in[9] = 1; act_sel_in[10] = 1; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 0; act_sel_in[14] = 0; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=5; act_sel_in[0] = 3; act_sel_in[1] = 2; act_sel_in[2] = 4; act_sel_in[3] = 2; act_sel_in[4] = 0; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 1; act_sel_in[8] = 0; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 1; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=4; act_sel_in[0] = 0; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 0; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 4; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=3; act_sel_in[0] = 3; act_sel_in[1] = 0; act_sel_in[2] = 0; act_sel_in[3] = 2; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 1; act_sel_in[11] = 4; act_sel_in[12] = 1; act_sel_in[13] = 2; act_sel_in[14] = 3; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=2; act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 3; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 1; act_sel_in[7] = 4; act_sel_in[8] = 4; act_sel_in[9] = 3; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=1; act_sel_in[0] = 2; act_sel_in[1] = 0; act_sel_in[2] = 4; act_sel_in[3] = 2; act_sel_in[4] = 2; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 3; act_sel_in[9] = 1; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 4; act_sel_in[13] = 4; act_sel_in[14] = 2; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 3; act_sel_in[1] = 2; act_sel_in[2] = 3; act_sel_in[3] = 2; act_sel_in[4] = 0; act_sel_in[5] = 0; act_sel_in[6] = 1; act_sel_in[7] = 3; act_sel_in[8] = 1; act_sel_in[9] = 0; act_sel_in[10] = 2; act_sel_in[11] = 1; act_sel_in[12] = 2; act_sel_in[13] = 2; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 


    #1 is_msb=1; column_idx=7; act_in[0] = 36; act_in[1] = 80; act_in[2] = 94; act_in[3] = -1; act_in[4] = 65; act_in[5] = 55; act_in[6] = -121; act_in[7] = 83; act_in[8] = -32; act_in[9] = 87; act_in[10] = -68; act_in[11] = 18; act_in[12] = 48; act_in[13] = 60; act_in[14] = -117; act_in[15] = -54; act_in[16] = -49; act_in[17] = 73; act_in[18] = -98; act_in[19] = 55; act_in[20] = 7; act_in[21] = -12; act_in[22] = 33; act_in[23] = 39; act_in[24] = -88; act_in[25] = -44; act_in[26] = 31; act_in[27] = 111; act_in[28] = -19; act_in[29] = -77; act_in[30] = -49; act_in[31] = 97; 
    act_sel_in[0] = 3; act_sel_in[1] = 1; act_sel_in[2] = 4; act_sel_in[3] = 3; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 4; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 1; act_sel_in[4] = 0; act_sel_in[5] = 1; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 3; act_sel_in[11] = 4; act_sel_in[12] = 1; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=5; act_sel_in[0] = 3; act_sel_in[1] = 0; act_sel_in[2] = 1; act_sel_in[3] = 3; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 4; act_sel_in[9] = 4; act_sel_in[10] = 4; act_sel_in[11] = 2; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=4; act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 2; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 0; act_sel_in[7] = 2; act_sel_in[8] = 1; act_sel_in[9] = 2; act_sel_in[10] = 0; act_sel_in[11] = 2; act_sel_in[12] = 0; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 2; act_sel_in[7] = 2; act_sel_in[8] = 3; act_sel_in[9] = 0; act_sel_in[10] = 4; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=2; act_sel_in[0] = 4; act_sel_in[1] = 4; act_sel_in[2] = 0; act_sel_in[3] = 3; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 4; act_sel_in[7] = 3; act_sel_in[8] = 1; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 4; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 3; act_sel_in[1] = 0; act_sel_in[2] = 0; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 3; act_sel_in[6] = 0; act_sel_in[7] = 3; act_sel_in[8] = 2; act_sel_in[9] = 0; act_sel_in[10] = 3; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 3; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=0; act_sel_in[0] = 2; act_sel_in[1] = 2; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 1; act_sel_in[5] = 4; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 3; act_sel_in[9] = 1; act_sel_in[10] = 4; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 4; act_sel_in[14] = 3; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 


    #1 is_msb=1; column_idx=7; act_in[0] = 40; act_in[1] = 9; act_in[2] = -86; act_in[3] = -10; act_in[4] = -43; act_in[5] = -55; act_in[6] = 64; act_in[7] = 17; act_in[8] = 70; act_in[9] = -75; act_in[10] = -90; act_in[11] = -94; act_in[12] = -67; act_in[13] = 89; act_in[14] = 86; act_in[15] = -104; act_in[16] = -26; act_in[17] = -23; act_in[18] = 50; act_in[19] = -117; act_in[20] = 118; act_in[21] = 72; act_in[22] = -124; act_in[23] = -79; act_in[24] = 50; act_in[25] = -96; act_in[26] = -80; act_in[27] = -125; act_in[28] = 55; act_in[29] = -71; act_in[30] = 2; act_in[31] = 104; 
    act_sel_in[0] = 4; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 2; act_sel_in[4] = 4; act_sel_in[5] = 1; act_sel_in[6] = 0; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 1; act_sel_in[14] = 3; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 0; act_sel_in[1] = 0; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 2; act_sel_in[5] = 4; act_sel_in[6] = 0; act_sel_in[7] = 4; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=5; act_sel_in[0] = 2; act_sel_in[1] = 0; act_sel_in[2] = 0; act_sel_in[3] = 1; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 1; act_sel_in[10] = 4; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 3; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=4; act_sel_in[0] = 3; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 3; act_sel_in[5] = 4; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 0; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 3; act_sel_in[1] = 2; act_sel_in[2] = 4; act_sel_in[3] = 3; act_sel_in[4] = 3; act_sel_in[5] = 1; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 4; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=2; act_sel_in[0] = 4; act_sel_in[1] = 0; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 0; act_sel_in[5] = 1; act_sel_in[6] = 0; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 4; act_sel_in[11] = 0; act_sel_in[12] = 4; act_sel_in[13] = 4; act_sel_in[14] = 3; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=1; act_sel_in[0] = 3; act_sel_in[1] = 0; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 3; act_sel_in[5] = 1; act_sel_in[6] = 3; act_sel_in[7] = 1; act_sel_in[8] = 3; act_sel_in[9] = 0; act_sel_in[10] = 3; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 1; act_sel_in[14] = 1; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 4; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 3; act_sel_in[8] = 3; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 1; act_sel_in[14] = 1; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 


    #1 is_msb=1; column_idx=7; act_in[0] = -105; act_in[1] = 91; act_in[2] = 92; act_in[3] = 35; act_in[4] = -32; act_in[5] = -7; act_in[6] = -2; act_in[7] = 48; act_in[8] = -59; act_in[9] = 13; act_in[10] = -89; act_in[11] = -91; act_in[12] = 108; act_in[13] = 35; act_in[14] = 93; act_in[15] = 0; act_in[16] = 21; act_in[17] = 97; act_in[18] = 115; act_in[19] = -93; act_in[20] = -100; act_in[21] = -98; act_in[22] = 111; act_in[23] = 111; act_in[24] = 8; act_in[25] = 81; act_in[26] = 30; act_in[27] = 80; act_in[28] = 74; act_in[29] = -39; act_in[30] = 86; act_in[31] = -73; 
    act_sel_in[0] = 3; act_sel_in[1] = 2; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 0; act_sel_in[5] = 0; act_sel_in[6] = 0; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 1; act_sel_in[10] = 1; act_sel_in[11] = 3; act_sel_in[12] = 1; act_sel_in[13] = 2; act_sel_in[14] = 3; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 2; act_sel_in[1] = 0; act_sel_in[2] = 4; act_sel_in[3] = 0; act_sel_in[4] = 4; act_sel_in[5] = 4; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 2; act_sel_in[9] = 4; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=5; act_sel_in[0] = 2; act_sel_in[1] = 3; act_sel_in[2] = 1; act_sel_in[3] = 3; act_sel_in[4] = 2; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 3; act_sel_in[8] = 4; act_sel_in[9] = 2; act_sel_in[10] = 2; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 3; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=4; act_sel_in[0] = 3; act_sel_in[1] = 0; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 3; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 2; act_sel_in[13] = 2; act_sel_in[14] = 1; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=3; act_sel_in[0] = 1; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 4; act_sel_in[4] = 1; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 1; act_sel_in[9] = 4; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 4; act_sel_in[14] = 1; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=2; act_sel_in[0] = 4; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 4; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 1; act_sel_in[9] = 2; act_sel_in[10] = 3; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 0; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=1; act_sel_in[0] = 4; act_sel_in[1] = 1; act_sel_in[2] = 4; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 3; act_sel_in[7] = 1; act_sel_in[8] = 2; act_sel_in[9] = 3; act_sel_in[10] = 1; act_sel_in[11] = 3; act_sel_in[12] = 0; act_sel_in[13] = 2; act_sel_in[14] = 1; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=0; act_sel_in[0] = 3; act_sel_in[1] = 2; act_sel_in[2] = 1; act_sel_in[3] = 4; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 3; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 


    #1 is_msb=1; column_idx=7; act_in[0] = -34; act_in[1] = 46; act_in[2] = -99; act_in[3] = 14; act_in[4] = 125; act_in[5] = -110; act_in[6] = -110; act_in[7] = -43; act_in[8] = -102; act_in[9] = 59; act_in[10] = -85; act_in[11] = 72; act_in[12] = 127; act_in[13] = 14; act_in[14] = -110; act_in[15] = -20; act_in[16] = 9; act_in[17] = -35; act_in[18] = -101; act_in[19] = -108; act_in[20] = -127; act_in[21] = 39; act_in[22] = -68; act_in[23] = 77; act_in[24] = 32; act_in[25] = -73; act_in[26] = -54; act_in[27] = -55; act_in[28] = 39; act_in[29] = -69; act_in[30] = 20; act_in[31] = 14; 
    act_sel_in[0] = 0; act_sel_in[1] = 0; act_sel_in[2] = 4; act_sel_in[3] = 0; act_sel_in[4] = 2; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 3; act_sel_in[8] = 2; act_sel_in[9] = 3; act_sel_in[10] = 0; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 4; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 2; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 2; act_sel_in[4] = 2; act_sel_in[5] = 1; act_sel_in[6] = 3; act_sel_in[7] = 1; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 4; act_sel_in[11] = 2; act_sel_in[12] = 3; act_sel_in[13] = 4; act_sel_in[14] = 1; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=5; act_sel_in[0] = 2; act_sel_in[1] = 0; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 1; act_sel_in[5] = 0; act_sel_in[6] = 1; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 0; act_sel_in[10] = 3; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 3; act_sel_in[14] = 3; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=4; act_sel_in[0] = 2; act_sel_in[1] = 0; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 3; act_sel_in[11] = 0; act_sel_in[12] = 1; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=3; act_sel_in[0] = 4; act_sel_in[1] = 3; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 2; act_sel_in[5] = 4; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 4; act_sel_in[12] = 4; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=2; act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 2; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 0; act_sel_in[6] = 0; act_sel_in[7] = 2; act_sel_in[8] = 3; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 3; act_sel_in[12] = 3; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 3; act_sel_in[1] = 0; act_sel_in[2] = 4; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 4; act_sel_in[11] = 2; act_sel_in[12] = 4; act_sel_in[13] = 1; act_sel_in[14] = 3; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=0; act_sel_in[0] = 4; act_sel_in[1] = 4; act_sel_in[2] = 4; act_sel_in[3] = 2; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 2; act_sel_in[7] = 3; act_sel_in[8] = 4; act_sel_in[9] = 0; act_sel_in[10] = 2; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 2; act_sel_in[14] = 1; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 


    #1 is_msb=1; column_idx=7; act_in[0] = -112; act_in[1] = 68; act_in[2] = -53; act_in[3] = 81; act_in[4] = 22; act_in[5] = -124; act_in[6] = 4; act_in[7] = 101; act_in[8] = 91; act_in[9] = -3; act_in[10] = -5; act_in[11] = -64; act_in[12] = -89; act_in[13] = -98; act_in[14] = -53; act_in[15] = 72; act_in[16] = 104; act_in[17] = 97; act_in[18] = -58; act_in[19] = 71; act_in[20] = -63; act_in[21] = 20; act_in[22] = 80; act_in[23] = 119; act_in[24] = 17; act_in[25] = -42; act_in[26] = 55; act_in[27] = -103; act_in[28] = 108; act_in[29] = -61; act_in[30] = -70; act_in[31] = -37; 
    act_sel_in[0] = 1; act_sel_in[1] = 0; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 4; act_sel_in[6] = 4; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 1; act_sel_in[11] = 3; act_sel_in[12] = 0; act_sel_in[13] = 2; act_sel_in[14] = 3; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 3; act_sel_in[1] = 0; act_sel_in[2] = 2; act_sel_in[3] = 1; act_sel_in[4] = 3; act_sel_in[5] = 0; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=5; act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 4; act_sel_in[3] = 0; act_sel_in[4] = 2; act_sel_in[5] = 4; act_sel_in[6] = 4; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 3; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 0; act_sel_in[14] = 1; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=4; act_sel_in[0] = 3; act_sel_in[1] = 3; act_sel_in[2] = 0; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 0; act_sel_in[7] = 2; act_sel_in[8] = 1; act_sel_in[9] = 2; act_sel_in[10] = 3; act_sel_in[11] = 2; act_sel_in[12] = 3; act_sel_in[13] = 4; act_sel_in[14] = 4; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 3; act_sel_in[1] = 3; act_sel_in[2] = 0; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 0; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 0; act_sel_in[10] = 2; act_sel_in[11] = 0; act_sel_in[12] = 3; act_sel_in[13] = 1; act_sel_in[14] = 3; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=2; act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 1; act_sel_in[6] = 1; act_sel_in[7] = 1; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 3; act_sel_in[11] = 4; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 1; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=1; act_sel_in[0] = 0; act_sel_in[1] = 0; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 1; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 3; act_sel_in[12] = 0; act_sel_in[13] = 2; act_sel_in[14] = 3; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 4; act_sel_in[1] = 4; act_sel_in[2] = 4; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 2; act_sel_in[7] = 3; act_sel_in[8] = 2; act_sel_in[9] = 3; act_sel_in[10] = 3; act_sel_in[11] = 0; act_sel_in[12] = 4; act_sel_in[13] = 4; act_sel_in[14] = 3; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 


    #1 is_msb=1; column_idx=7; act_in[0] = 64; act_in[1] = -43; act_in[2] = 77; act_in[3] = 62; act_in[4] = -20; act_in[5] = 84; act_in[6] = 16; act_in[7] = -119; act_in[8] = 73; act_in[9] = -107; act_in[10] = -39; act_in[11] = 16; act_in[12] = 27; act_in[13] = -102; act_in[14] = 24; act_in[15] = 0; act_in[16] = 56; act_in[17] = 5; act_in[18] = 125; act_in[19] = -106; act_in[20] = 90; act_in[21] = -126; act_in[22] = 49; act_in[23] = 44; act_in[24] = 10; act_in[25] = 77; act_in[26] = -104; act_in[27] = -86; act_in[28] = -52; act_in[29] = -54; act_in[30] = -73; act_in[31] = -5; 
    act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 4; act_sel_in[11] = 3; act_sel_in[12] = 4; act_sel_in[13] = 1; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 3; act_sel_in[1] = 3; act_sel_in[2] = 1; act_sel_in[3] = 3; act_sel_in[4] = 3; act_sel_in[5] = 0; act_sel_in[6] = 1; act_sel_in[7] = 3; act_sel_in[8] = 4; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 0; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=5; act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 1; act_sel_in[9] = 0; act_sel_in[10] = 2; act_sel_in[11] = 2; act_sel_in[12] = 3; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=4; act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 1; act_sel_in[9] = 2; act_sel_in[10] = 0; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 0; act_sel_in[14] = 1; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=3; act_sel_in[0] = 3; act_sel_in[1] = 2; act_sel_in[2] = 1; act_sel_in[3] = 0; act_sel_in[4] = 2; act_sel_in[5] = 1; act_sel_in[6] = 1; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 1; act_sel_in[11] = 0; act_sel_in[12] = 3; act_sel_in[13] = 4; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=2; act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 3; act_sel_in[3] = 2; act_sel_in[4] = 4; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 4; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 3; act_sel_in[11] = 2; act_sel_in[12] = 3; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 1; act_sel_in[1] = 0; act_sel_in[2] = 2; act_sel_in[3] = 2; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 4; act_sel_in[7] = 3; act_sel_in[8] = 4; act_sel_in[9] = 0; act_sel_in[10] = 0; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 1; act_sel_in[14] = 3; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 3; act_sel_in[1] = 0; act_sel_in[2] = 1; act_sel_in[3] = 0; act_sel_in[4] = 0; act_sel_in[5] = 2; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 1; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 2; act_sel_in[14] = 3; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 


    #1 is_msb=1; column_idx=7; act_in[0] = -23; act_in[1] = -20; act_in[2] = 125; act_in[3] = 4; act_in[4] = 119; act_in[5] = -104; act_in[6] = 79; act_in[7] = -45; act_in[8] = 118; act_in[9] = -6; act_in[10] = -84; act_in[11] = 73; act_in[12] = -105; act_in[13] = -104; act_in[14] = -71; act_in[15] = -36; act_in[16] = 70; act_in[17] = 81; act_in[18] = 54; act_in[19] = 45; act_in[20] = -25; act_in[21] = -86; act_in[22] = -47; act_in[23] = 2; act_in[24] = -13; act_in[25] = 31; act_in[26] = -81; act_in[27] = -42; act_in[28] = 56; act_in[29] = -57; act_in[30] = -67; act_in[31] = -44; 
    act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 0; act_sel_in[11] = 2; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 3; act_sel_in[1] = 4; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 2; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 4; act_sel_in[12] = 1; act_sel_in[13] = 0; act_sel_in[14] = 3; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=5; act_sel_in[0] = 1; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 3; act_sel_in[8] = 2; act_sel_in[9] = 0; act_sel_in[10] = 3; act_sel_in[11] = 3; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 1; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=4; act_sel_in[0] = 3; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 2; act_sel_in[4] = 0; act_sel_in[5] = 2; act_sel_in[6] = 0; act_sel_in[7] = 0; act_sel_in[8] = 3; act_sel_in[9] = 0; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 3; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=3; act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 2; act_sel_in[3] = 0; act_sel_in[4] = 4; act_sel_in[5] = 4; act_sel_in[6] = 2; act_sel_in[7] = 4; act_sel_in[8] = 4; act_sel_in[9] = 0; act_sel_in[10] = 3; act_sel_in[11] = 4; act_sel_in[12] = 4; act_sel_in[13] = 3; act_sel_in[14] = 3; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=2; act_sel_in[0] = 4; act_sel_in[1] = 3; act_sel_in[2] = 4; act_sel_in[3] = 2; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 1; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 4; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=1; act_sel_in[0] = 2; act_sel_in[1] = 0; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 1; act_sel_in[5] = 4; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 2; act_sel_in[9] = 1; act_sel_in[10] = 3; act_sel_in[11] = 2; act_sel_in[12] = 3; act_sel_in[13] = 1; act_sel_in[14] = 3; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 3; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 1; act_sel_in[11] = 3; act_sel_in[12] = 4; act_sel_in[13] = 4; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 


    #1 is_msb=1; column_idx=7; act_in[0] = -5; act_in[1] = 47; act_in[2] = 9; act_in[3] = 19; act_in[4] = -106; act_in[5] = -120; act_in[6] = 64; act_in[7] = -113; act_in[8] = -1; act_in[9] = -71; act_in[10] = -61; act_in[11] = -55; act_in[12] = 113; act_in[13] = 87; act_in[14] = -31; act_in[15] = -67; act_in[16] = 79; act_in[17] = 35; act_in[18] = 30; act_in[19] = 90; act_in[20] = -34; act_in[21] = -17; act_in[22] = -71; act_in[23] = 64; act_in[24] = 56; act_in[25] = 101; act_in[26] = -75; act_in[27] = -119; act_in[28] = -100; act_in[29] = 49; act_in[30] = -128; act_in[31] = -10; 
    act_sel_in[0] = 2; act_sel_in[1] = 4; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 4; act_sel_in[6] = 4; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 1; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 1; act_sel_in[1] = 1; act_sel_in[2] = 4; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 1; act_sel_in[6] = 1; act_sel_in[7] = 4; act_sel_in[8] = 1; act_sel_in[9] = 1; act_sel_in[10] = 4; act_sel_in[11] = 3; act_sel_in[12] = 2; act_sel_in[13] = 0; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=5; act_sel_in[0] = 1; act_sel_in[1] = 4; act_sel_in[2] = 1; act_sel_in[3] = 3; act_sel_in[4] = 0; act_sel_in[5] = 1; act_sel_in[6] = 3; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 2; act_sel_in[11] = 4; act_sel_in[12] = 3; act_sel_in[13] = 0; act_sel_in[14] = 4; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=4; act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 2; act_sel_in[6] = 3; act_sel_in[7] = 1; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 2; act_sel_in[14] = 0; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=3; act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 0; act_sel_in[3] = 0; act_sel_in[4] = 2; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 3; act_sel_in[11] = 0; act_sel_in[12] = 3; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=2; act_sel_in[0] = 4; act_sel_in[1] = 3; act_sel_in[2] = 1; act_sel_in[3] = 4; act_sel_in[4] = 0; act_sel_in[5] = 4; act_sel_in[6] = 1; act_sel_in[7] = 1; act_sel_in[8] = 4; act_sel_in[9] = 4; act_sel_in[10] = 3; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 2; act_sel_in[14] = 1; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 4; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 4; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 1; act_sel_in[14] = 0; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 1; act_sel_in[4] = 0; act_sel_in[5] = 1; act_sel_in[6] = 1; act_sel_in[7] = 4; act_sel_in[8] = 2; act_sel_in[9] = 3; act_sel_in[10] = 1; act_sel_in[11] = 0; act_sel_in[12] = 3; act_sel_in[13] = 4; act_sel_in[14] = 1; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 


    #1 is_msb=1; column_idx=7; act_in[0] = -22; act_in[1] = -13; act_in[2] = 20; act_in[3] = 15; act_in[4] = -21; act_in[5] = 36; act_in[6] = 115; act_in[7] = 52; act_in[8] = -59; act_in[9] = 67; act_in[10] = -80; act_in[11] = -39; act_in[12] = 101; act_in[13] = 29; act_in[14] = -44; act_in[15] = -10; act_in[16] = 81; act_in[17] = -19; act_in[18] = -86; act_in[19] = -57; act_in[20] = -52; act_in[21] = 55; act_in[22] = -69; act_in[23] = 89; act_in[24] = 7; act_in[25] = -117; act_in[26] = 1; act_in[27] = 92; act_in[28] = 10; act_in[29] = 48; act_in[30] = -104; act_in[31] = -44; 
    act_sel_in[0] = 3; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 4; act_sel_in[6] = 2; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 1; act_sel_in[10] = 4; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 1; act_sel_in[14] = 1; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 3; act_sel_in[1] = 1; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 3; act_sel_in[10] = 1; act_sel_in[11] = 1; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=5; act_sel_in[0] = 0; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 3; act_sel_in[10] = 2; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 3; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=4; act_sel_in[0] = 4; act_sel_in[1] = 1; act_sel_in[2] = 0; act_sel_in[3] = 0; act_sel_in[4] = 0; act_sel_in[5] = 3; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 4; act_sel_in[9] = 0; act_sel_in[10] = 3; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 4; act_sel_in[14] = 1; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 4; act_sel_in[5] = 4; act_sel_in[6] = 1; act_sel_in[7] = 1; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 4; act_sel_in[14] = 4; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=2; act_sel_in[0] = 3; act_sel_in[1] = 3; act_sel_in[2] = 0; act_sel_in[3] = 0; act_sel_in[4] = 4; act_sel_in[5] = 4; act_sel_in[6] = 2; act_sel_in[7] = 2; act_sel_in[8] = 4; act_sel_in[9] = 4; act_sel_in[10] = 0; act_sel_in[11] = 4; act_sel_in[12] = 4; act_sel_in[13] = 3; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=1; act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 1; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 0; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 3; act_sel_in[11] = 4; act_sel_in[12] = 1; act_sel_in[13] = 4; act_sel_in[14] = 2; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=0; act_sel_in[0] = 4; act_sel_in[1] = 0; act_sel_in[2] = 4; act_sel_in[3] = 1; act_sel_in[4] = 3; act_sel_in[5] = 1; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 3; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 2; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 


    #1 is_msb=1; column_idx=7; act_in[0] = 83; act_in[1] = 64; act_in[2] = -90; act_in[3] = -20; act_in[4] = -24; act_in[5] = 92; act_in[6] = 43; act_in[7] = 15; act_in[8] = 91; act_in[9] = -60; act_in[10] = 2; act_in[11] = -75; act_in[12] = 125; act_in[13] = -125; act_in[14] = 52; act_in[15] = -2; act_in[16] = 21; act_in[17] = -71; act_in[18] = 50; act_in[19] = -63; act_in[20] = -23; act_in[21] = -19; act_in[22] = -25; act_in[23] = -48; act_in[24] = 71; act_in[25] = -91; act_in[26] = -81; act_in[27] = 121; act_in[28] = -120; act_in[29] = 118; act_in[30] = 37; act_in[31] = 82; 
    act_sel_in[0] = 3; act_sel_in[1] = 2; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 2; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 1; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 0; act_sel_in[13] = 2; act_sel_in[14] = 1; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 1; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 2; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 2; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 2; act_sel_in[12] = 0; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=5; act_sel_in[0] = 1; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 0; act_sel_in[5] = 2; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 2; act_sel_in[14] = 3; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=4; act_sel_in[0] = 4; act_sel_in[1] = 0; act_sel_in[2] = 3; act_sel_in[3] = 4; act_sel_in[4] = 0; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 4; act_sel_in[9] = 3; act_sel_in[10] = 0; act_sel_in[11] = 3; act_sel_in[12] = 3; act_sel_in[13] = 0; act_sel_in[14] = 1; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 3; act_sel_in[1] = 3; act_sel_in[2] = 0; act_sel_in[3] = 1; act_sel_in[4] = 0; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 3; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 0; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=2; act_sel_in[0] = 2; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 2; act_sel_in[4] = 0; act_sel_in[5] = 4; act_sel_in[6] = 0; act_sel_in[7] = 1; act_sel_in[8] = 1; act_sel_in[9] = 3; act_sel_in[10] = 1; act_sel_in[11] = 3; act_sel_in[12] = 2; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 0; act_sel_in[3] = 3; act_sel_in[4] = 4; act_sel_in[5] = 4; act_sel_in[6] = 4; act_sel_in[7] = 3; act_sel_in[8] = 2; act_sel_in[9] = 0; act_sel_in[10] = 0; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 4; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 4; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 0; act_sel_in[7] = 1; act_sel_in[8] = 1; act_sel_in[9] = 0; act_sel_in[10] = 2; act_sel_in[11] = 3; act_sel_in[12] = 0; act_sel_in[13] = 2; act_sel_in[14] = 3; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 


    #1 is_msb=1; column_idx=7; act_in[0] = 92; act_in[1] = -119; act_in[2] = -71; act_in[3] = -119; act_in[4] = 62; act_in[5] = 3; act_in[6] = -14; act_in[7] = -45; act_in[8] = 113; act_in[9] = 77; act_in[10] = 13; act_in[11] = -12; act_in[12] = -52; act_in[13] = -6; act_in[14] = -31; act_in[15] = -53; act_in[16] = 113; act_in[17] = 66; act_in[18] = 44; act_in[19] = 3; act_in[20] = -74; act_in[21] = -62; act_in[22] = -6; act_in[23] = -15; act_in[24] = -47; act_in[25] = -56; act_in[26] = -6; act_in[27] = 84; act_in[28] = -71; act_in[29] = 48; act_in[30] = -71; act_in[31] = 24; 
    act_sel_in[0] = 4; act_sel_in[1] = 0; act_sel_in[2] = 3; act_sel_in[3] = 2; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 1; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 3; act_sel_in[11] = 0; act_sel_in[12] = 1; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 3; act_sel_in[1] = 2; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 2; act_sel_in[7] = 4; act_sel_in[8] = 1; act_sel_in[9] = 3; act_sel_in[10] = 3; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 1; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=5; act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 3; act_sel_in[3] = 2; act_sel_in[4] = 2; act_sel_in[5] = 3; act_sel_in[6] = 0; act_sel_in[7] = 4; act_sel_in[8] = 1; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 1; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=4; act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 2; act_sel_in[3] = 3; act_sel_in[4] = 3; act_sel_in[5] = 0; act_sel_in[6] = 0; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 2; act_sel_in[10] = 3; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 1; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 2; act_sel_in[4] = 0; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 4; act_sel_in[11] = 3; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=2; act_sel_in[0] = 2; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 2; act_sel_in[4] = 3; act_sel_in[5] = 4; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 3; act_sel_in[10] = 0; act_sel_in[11] = 2; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 2; act_sel_in[1] = 4; act_sel_in[2] = 4; act_sel_in[3] = 0; act_sel_in[4] = 0; act_sel_in[5] = 4; act_sel_in[6] = 0; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 2; act_sel_in[11] = 0; act_sel_in[12] = 4; act_sel_in[13] = 3; act_sel_in[14] = 0; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 2; act_sel_in[3] = 0; act_sel_in[4] = 4; act_sel_in[5] = 1; act_sel_in[6] = 0; act_sel_in[7] = 4; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 4; act_sel_in[14] = 3; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 


    #1 is_msb=1; column_idx=7; act_in[0] = 22; act_in[1] = 47; act_in[2] = 62; act_in[3] = 9; act_in[4] = 96; act_in[5] = -73; act_in[6] = 80; act_in[7] = -24; act_in[8] = -34; act_in[9] = 113; act_in[10] = -73; act_in[11] = 25; act_in[12] = -66; act_in[13] = 95; act_in[14] = 50; act_in[15] = -49; act_in[16] = 38; act_in[17] = -89; act_in[18] = 101; act_in[19] = -42; act_in[20] = -27; act_in[21] = 75; act_in[22] = 44; act_in[23] = -17; act_in[24] = 24; act_in[25] = 44; act_in[26] = 77; act_in[27] = 104; act_in[28] = -96; act_in[29] = 57; act_in[30] = 69; act_in[31] = 90; 
    act_sel_in[0] = 0; act_sel_in[1] = 1; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 2; act_sel_in[5] = 3; act_sel_in[6] = 2; act_sel_in[7] = 2; act_sel_in[8] = 4; act_sel_in[9] = 4; act_sel_in[10] = 4; act_sel_in[11] = 4; act_sel_in[12] = 1; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 0; act_sel_in[1] = 0; act_sel_in[2] = 0; act_sel_in[3] = 2; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 4; act_sel_in[9] = 0; act_sel_in[10] = 2; act_sel_in[11] = 0; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 3; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=5; act_sel_in[0] = 4; act_sel_in[1] = 0; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 1; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 0; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 0; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=4; act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 4; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 3; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 0; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 1; act_sel_in[1] = 1; act_sel_in[2] = 0; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 2; act_sel_in[8] = 3; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=2; act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 0; act_sel_in[3] = 1; act_sel_in[4] = 3; act_sel_in[5] = 1; act_sel_in[6] = 2; act_sel_in[7] = 3; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 3; act_sel_in[11] = 3; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 3; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 0; act_sel_in[12] = 4; act_sel_in[13] = 0; act_sel_in[14] = 3; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 1; act_sel_in[5] = 4; act_sel_in[6] = 1; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 3; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 4; act_sel_in[14] = 3; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 


    #1 is_msb=1; column_idx=7; act_in[0] = -53; act_in[1] = 125; act_in[2] = 118; act_in[3] = -118; act_in[4] = 71; act_in[5] = -3; act_in[6] = 16; act_in[7] = -31; act_in[8] = -17; act_in[9] = 3; act_in[10] = 93; act_in[11] = 58; act_in[12] = -14; act_in[13] = -97; act_in[14] = 120; act_in[15] = -18; act_in[16] = -113; act_in[17] = 49; act_in[18] = 103; act_in[19] = -102; act_in[20] = 0; act_in[21] = 18; act_in[22] = 19; act_in[23] = 1; act_in[24] = -6; act_in[25] = 10; act_in[26] = -39; act_in[27] = -32; act_in[28] = -50; act_in[29] = 83; act_in[30] = 30; act_in[31] = -75; 
    act_sel_in[0] = 4; act_sel_in[1] = 3; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 4; act_sel_in[6] = 4; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 3; act_sel_in[12] = 0; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 2; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 3; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 3; act_sel_in[12] = 2; act_sel_in[13] = 2; act_sel_in[14] = 3; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=5; act_sel_in[0] = 3; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 4; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 2; act_sel_in[13] = 1; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=4; act_sel_in[0] = 2; act_sel_in[1] = 0; act_sel_in[2] = 2; act_sel_in[3] = 2; act_sel_in[4] = 2; act_sel_in[5] = 4; act_sel_in[6] = 1; act_sel_in[7] = 1; act_sel_in[8] = 1; act_sel_in[9] = 1; act_sel_in[10] = 4; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=3; act_sel_in[0] = 1; act_sel_in[1] = 4; act_sel_in[2] = 0; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 1; act_sel_in[6] = 1; act_sel_in[7] = 3; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 2; act_sel_in[12] = 3; act_sel_in[13] = 4; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=2; act_sel_in[0] = 4; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 4; act_sel_in[6] = 1; act_sel_in[7] = 3; act_sel_in[8] = 4; act_sel_in[9] = 0; act_sel_in[10] = 0; act_sel_in[11] = 4; act_sel_in[12] = 4; act_sel_in[13] = 0; act_sel_in[14] = 3; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 3; act_sel_in[1] = 2; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 1; act_sel_in[8] = 1; act_sel_in[9] = 2; act_sel_in[10] = 0; act_sel_in[11] = 0; act_sel_in[12] = 1; act_sel_in[13] = 0; act_sel_in[14] = 0; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 3; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 3; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 1; act_sel_in[7] = 3; act_sel_in[8] = 4; act_sel_in[9] = 3; act_sel_in[10] = 0; act_sel_in[11] = 2; act_sel_in[12] = 3; act_sel_in[13] = 2; act_sel_in[14] = 3; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 


    #1 is_msb=1; column_idx=7; act_in[0] = 94; act_in[1] = 105; act_in[2] = 89; act_in[3] = 127; act_in[4] = -116; act_in[5] = 53; act_in[6] = -53; act_in[7] = 28; act_in[8] = -47; act_in[9] = -65; act_in[10] = -33; act_in[11] = 32; act_in[12] = 15; act_in[13] = -44; act_in[14] = -77; act_in[15] = -7; act_in[16] = 54; act_in[17] = -22; act_in[18] = 19; act_in[19] = 41; act_in[20] = -60; act_in[21] = -119; act_in[22] = -66; act_in[23] = -57; act_in[24] = 3; act_in[25] = -30; act_in[26] = -35; act_in[27] = -48; act_in[28] = -123; act_in[29] = -16; act_in[30] = -82; act_in[31] = 14; 
    act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 3; act_sel_in[3] = 2; act_sel_in[4] = 3; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 2; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 1; act_sel_in[11] = 1; act_sel_in[12] = 2; act_sel_in[13] = 1; act_sel_in[14] = 1; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 1; act_sel_in[3] = 4; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 3; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 4; act_sel_in[14] = 3; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=5; act_sel_in[0] = 0; act_sel_in[1] = 0; act_sel_in[2] = 4; act_sel_in[3] = 1; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 1; act_sel_in[7] = 1; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 3; act_sel_in[11] = 0; act_sel_in[12] = 3; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=4; act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 0; act_sel_in[5] = 1; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 2; act_sel_in[9] = 4; act_sel_in[10] = 0; act_sel_in[11] = 2; act_sel_in[12] = 3; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=3; act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 4; act_sel_in[6] = 0; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 3; act_sel_in[12] = 0; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=2; act_sel_in[0] = 2; act_sel_in[1] = 0; act_sel_in[2] = 1; act_sel_in[3] = 4; act_sel_in[4] = 2; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 2; act_sel_in[8] = 4; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 1; act_sel_in[12] = 2; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 0; act_sel_in[7] = 3; act_sel_in[8] = 1; act_sel_in[9] = 3; act_sel_in[10] = 1; act_sel_in[11] = 3; act_sel_in[12] = 3; act_sel_in[13] = 0; act_sel_in[14] = 3; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 1; act_sel_in[1] = 4; act_sel_in[2] = 4; act_sel_in[3] = 2; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 2; act_sel_in[10] = 2; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 


    #1 is_msb=1; column_idx=7; act_in[0] = 108; act_in[1] = 122; act_in[2] = 25; act_in[3] = 31; act_in[4] = -84; act_in[5] = -84; act_in[6] = 48; act_in[7] = -102; act_in[8] = 33; act_in[9] = -43; act_in[10] = -109; act_in[11] = 39; act_in[12] = -18; act_in[13] = 127; act_in[14] = -122; act_in[15] = -72; act_in[16] = 45; act_in[17] = 72; act_in[18] = -11; act_in[19] = 121; act_in[20] = -35; act_in[21] = 91; act_in[22] = -122; act_in[23] = -29; act_in[24] = -121; act_in[25] = -48; act_in[26] = -127; act_in[27] = 125; act_in[28] = -103; act_in[29] = -58; act_in[30] = -8; act_in[31] = 115; 
    act_sel_in[0] = 1; act_sel_in[1] = 0; act_sel_in[2] = 2; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 4; act_sel_in[9] = 3; act_sel_in[10] = 1; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 4; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 3; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 0; act_sel_in[7] = 2; act_sel_in[8] = 1; act_sel_in[9] = 3; act_sel_in[10] = 2; act_sel_in[11] = 4; act_sel_in[12] = 1; act_sel_in[13] = 0; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=5; act_sel_in[0] = 2; act_sel_in[1] = 0; act_sel_in[2] = 4; act_sel_in[3] = 3; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 0; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 1; act_sel_in[14] = 3; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=4; act_sel_in[0] = 3; act_sel_in[1] = 3; act_sel_in[2] = 4; act_sel_in[3] = 2; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 4; act_sel_in[7] = 3; act_sel_in[8] = 2; act_sel_in[9] = 0; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 0; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 1; act_sel_in[3] = 4; act_sel_in[4] = 2; act_sel_in[5] = 2; act_sel_in[6] = 3; act_sel_in[7] = 2; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 3; act_sel_in[12] = 3; act_sel_in[13] = 3; act_sel_in[14] = 3; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=2; act_sel_in[0] = 4; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 0; act_sel_in[4] = 0; act_sel_in[5] = 0; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 2; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 0; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=1; act_sel_in[0] = 0; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 0; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 3; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 0; act_sel_in[1] = 1; act_sel_in[2] = 4; act_sel_in[3] = 2; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 2; act_sel_in[9] = 1; act_sel_in[10] = 3; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 


    #1 is_msb=1; column_idx=7; act_in[0] = 104; act_in[1] = 90; act_in[2] = 106; act_in[3] = -15; act_in[4] = -125; act_in[5] = 88; act_in[6] = 82; act_in[7] = -123; act_in[8] = 80; act_in[9] = 66; act_in[10] = 21; act_in[11] = -6; act_in[12] = 41; act_in[13] = -118; act_in[14] = 46; act_in[15] = -4; act_in[16] = -45; act_in[17] = -101; act_in[18] = 104; act_in[19] = -33; act_in[20] = -99; act_in[21] = -69; act_in[22] = 96; act_in[23] = -22; act_in[24] = 20; act_in[25] = -88; act_in[26] = -32; act_in[27] = -120; act_in[28] = -14; act_in[29] = 7; act_in[30] = 10; act_in[31] = 112; 
    act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 4; act_sel_in[3] = 0; act_sel_in[4] = 0; act_sel_in[5] = 1; act_sel_in[6] = 0; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 1; act_sel_in[12] = 2; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 2; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 2; act_sel_in[11] = 0; act_sel_in[12] = 3; act_sel_in[13] = 3; act_sel_in[14] = 3; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=5; act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 1; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 3; act_sel_in[9] = 0; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 0; act_sel_in[14] = 3; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=4; act_sel_in[0] = 3; act_sel_in[1] = 0; act_sel_in[2] = 2; act_sel_in[3] = 2; act_sel_in[4] = 2; act_sel_in[5] = 4; act_sel_in[6] = 1; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 2; act_sel_in[1] = 2; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 3; act_sel_in[9] = 1; act_sel_in[10] = 4; act_sel_in[11] = 3; act_sel_in[12] = 1; act_sel_in[13] = 4; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=2; act_sel_in[0] = 0; act_sel_in[1] = 0; act_sel_in[2] = 0; act_sel_in[3] = 0; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 2; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 3; act_sel_in[12] = 4; act_sel_in[13] = 3; act_sel_in[14] = 1; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 3; act_sel_in[3] = 2; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 3; act_sel_in[7] = 1; act_sel_in[8] = 1; act_sel_in[9] = 0; act_sel_in[10] = 3; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 0; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=0; act_sel_in[0] = 2; act_sel_in[1] = 0; act_sel_in[2] = 1; act_sel_in[3] = 3; act_sel_in[4] = 2; act_sel_in[5] = 0; act_sel_in[6] = 0; act_sel_in[7] = 1; act_sel_in[8] = 1; act_sel_in[9] = 0; act_sel_in[10] = 1; act_sel_in[11] = 1; act_sel_in[12] = 0; act_sel_in[13] = 0; act_sel_in[14] = 0; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 


    #1 is_msb=1; column_idx=7; act_in[0] = -120; act_in[1] = 10; act_in[2] = -113; act_in[3] = 69; act_in[4] = 84; act_in[5] = 98; act_in[6] = 14; act_in[7] = -48; act_in[8] = -91; act_in[9] = -58; act_in[10] = -100; act_in[11] = 29; act_in[12] = -115; act_in[13] = 12; act_in[14] = 7; act_in[15] = -39; act_in[16] = 107; act_in[17] = -57; act_in[18] = -105; act_in[19] = -101; act_in[20] = -72; act_in[21] = -23; act_in[22] = 59; act_in[23] = -38; act_in[24] = -78; act_in[25] = -17; act_in[26] = 35; act_in[27] = 93; act_in[28] = 104; act_in[29] = -14; act_in[30] = 31; act_in[31] = -128; 
    act_sel_in[0] = 1; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 2; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 0; act_sel_in[7] = 3; act_sel_in[8] = 1; act_sel_in[9] = 4; act_sel_in[10] = 0; act_sel_in[11] = 4; act_sel_in[12] = 1; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 0; act_sel_in[3] = 3; act_sel_in[4] = 2; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 4; act_sel_in[9] = 3; act_sel_in[10] = 0; act_sel_in[11] = 3; act_sel_in[12] = 4; act_sel_in[13] = 4; act_sel_in[14] = 3; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=5; act_sel_in[0] = 1; act_sel_in[1] = 0; act_sel_in[2] = 4; act_sel_in[3] = 3; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 3; act_sel_in[7] = 1; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 1; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 3; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=4; act_sel_in[0] = 4; act_sel_in[1] = 4; act_sel_in[2] = 4; act_sel_in[3] = 4; act_sel_in[4] = 0; act_sel_in[5] = 3; act_sel_in[6] = 4; act_sel_in[7] = 4; act_sel_in[8] = 1; act_sel_in[9] = 1; act_sel_in[10] = 3; act_sel_in[11] = 3; act_sel_in[12] = 4; act_sel_in[13] = 0; act_sel_in[14] = 3; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=3; act_sel_in[0] = 0; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 4; act_sel_in[12] = 3; act_sel_in[13] = 1; act_sel_in[14] = 1; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=2; act_sel_in[0] = 2; act_sel_in[1] = 0; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 0; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 2; act_sel_in[8] = 3; act_sel_in[9] = 2; act_sel_in[10] = 2; act_sel_in[11] = 2; act_sel_in[12] = 3; act_sel_in[13] = 3; act_sel_in[14] = 1; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 1; act_sel_in[1] = 0; act_sel_in[2] = 4; act_sel_in[3] = 3; act_sel_in[4] = 2; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 3; act_sel_in[8] = 4; act_sel_in[9] = 4; act_sel_in[10] = 4; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 2; act_sel_in[3] = 3; act_sel_in[4] = 1; act_sel_in[5] = 4; act_sel_in[6] = 0; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 2; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 


    #1 is_msb=1; column_idx=7; act_in[0] = 105; act_in[1] = -50; act_in[2] = 121; act_in[3] = 47; act_in[4] = -98; act_in[5] = -20; act_in[6] = 113; act_in[7] = 23; act_in[8] = -120; act_in[9] = 89; act_in[10] = 21; act_in[11] = -64; act_in[12] = -115; act_in[13] = 6; act_in[14] = 35; act_in[15] = -11; act_in[16] = -122; act_in[17] = 127; act_in[18] = 12; act_in[19] = 85; act_in[20] = -95; act_in[21] = -88; act_in[22] = 92; act_in[23] = -101; act_in[24] = -71; act_in[25] = 90; act_in[26] = 83; act_in[27] = 120; act_in[28] = 97; act_in[29] = 52; act_in[30] = -68; act_in[31] = -67; 
    act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 3; act_sel_in[8] = 1; act_sel_in[9] = 1; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 0; act_sel_in[1] = 1; act_sel_in[2] = 2; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 1; act_sel_in[6] = 1; act_sel_in[7] = 3; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 2; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=5; act_sel_in[0] = 0; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 2; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 3; act_sel_in[11] = 0; act_sel_in[12] = 3; act_sel_in[13] = 4; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=4; act_sel_in[0] = 3; act_sel_in[1] = 0; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 0; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 1; act_sel_in[11] = 4; act_sel_in[12] = 1; act_sel_in[13] = 3; act_sel_in[14] = 3; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 4; act_sel_in[1] = 0; act_sel_in[2] = 1; act_sel_in[3] = 3; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 0; act_sel_in[7] = 4; act_sel_in[8] = 2; act_sel_in[9] = 3; act_sel_in[10] = 1; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 0; act_sel_in[14] = 1; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=2; act_sel_in[0] = 3; act_sel_in[1] = 4; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 2; act_sel_in[5] = 3; act_sel_in[6] = 4; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 3; act_sel_in[11] = 3; act_sel_in[12] = 3; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 2; act_sel_in[1] = 2; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 0; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 4; act_sel_in[9] = 0; act_sel_in[10] = 4; act_sel_in[11] = 0; act_sel_in[12] = 3; act_sel_in[13] = 1; act_sel_in[14] = 0; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=0; act_sel_in[0] = 0; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 4; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 2; act_sel_in[11] = 1; act_sel_in[12] = 2; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 


    #1 is_msb=1; column_idx=7; act_in[0] = 31; act_in[1] = -6; act_in[2] = -112; act_in[3] = 5; act_in[4] = -124; act_in[5] = 32; act_in[6] = 50; act_in[7] = 95; act_in[8] = 120; act_in[9] = 2; act_in[10] = -81; act_in[11] = 115; act_in[12] = -6; act_in[13] = -42; act_in[14] = -105; act_in[15] = 120; act_in[16] = 3; act_in[17] = -10; act_in[18] = -2; act_in[19] = -89; act_in[20] = -64; act_in[21] = 96; act_in[22] = 84; act_in[23] = 121; act_in[24] = -16; act_in[25] = 109; act_in[26] = 57; act_in[27] = 58; act_in[28] = 70; act_in[29] = 34; act_in[30] = 25; act_in[31] = -84; 
    act_sel_in[0] = 1; act_sel_in[1] = 4; act_sel_in[2] = 0; act_sel_in[3] = 0; act_sel_in[4] = 0; act_sel_in[5] = 3; act_sel_in[6] = 2; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 2; act_sel_in[11] = 4; act_sel_in[12] = 3; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 4; act_sel_in[1] = 1; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 4; act_sel_in[9] = 3; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=5; act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 2; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 0; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 1; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 4; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=4; act_sel_in[0] = 2; act_sel_in[1] = 3; act_sel_in[2] = 4; act_sel_in[3] = 1; act_sel_in[4] = 1; act_sel_in[5] = 0; act_sel_in[6] = 4; act_sel_in[7] = 0; act_sel_in[8] = 4; act_sel_in[9] = 0; act_sel_in[10] = 0; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 0; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=3; act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 2; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 2; act_sel_in[9] = 0; act_sel_in[10] = 3; act_sel_in[11] = 0; act_sel_in[12] = 3; act_sel_in[13] = 0; act_sel_in[14] = 3; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=2; act_sel_in[0] = 4; act_sel_in[1] = 1; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 0; act_sel_in[5] = 4; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 3; act_sel_in[11] = 4; act_sel_in[12] = 1; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 1; act_sel_in[7] = 4; act_sel_in[8] = 4; act_sel_in[9] = 2; act_sel_in[10] = 2; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 3; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 1; act_sel_in[3] = 0; act_sel_in[4] = 4; act_sel_in[5] = 1; act_sel_in[6] = 0; act_sel_in[7] = 1; act_sel_in[8] = 3; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 0; act_sel_in[12] = 4; act_sel_in[13] = 0; act_sel_in[14] = 3; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 


    #1 is_msb=1; column_idx=7; act_in[0] = -89; act_in[1] = -90; act_in[2] = -105; act_in[3] = -87; act_in[4] = 9; act_in[5] = 40; act_in[6] = -114; act_in[7] = 0; act_in[8] = 125; act_in[9] = -98; act_in[10] = -21; act_in[11] = -19; act_in[12] = -7; act_in[13] = -124; act_in[14] = 7; act_in[15] = 117; act_in[16] = 59; act_in[17] = 61; act_in[18] = 9; act_in[19] = -3; act_in[20] = 81; act_in[21] = -122; act_in[22] = -115; act_in[23] = -4; act_in[24] = 87; act_in[25] = 43; act_in[26] = -45; act_in[27] = 43; act_in[28] = 80; act_in[29] = 80; act_in[30] = 13; act_in[31] = 105; 
    act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 0; act_sel_in[5] = 4; act_sel_in[6] = 2; act_sel_in[7] = 2; act_sel_in[8] = 0; act_sel_in[9] = 4; act_sel_in[10] = 3; act_sel_in[11] = 4; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 1; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 3; act_sel_in[8] = 2; act_sel_in[9] = 4; act_sel_in[10] = 0; act_sel_in[11] = 2; act_sel_in[12] = 4; act_sel_in[13] = 4; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=5; act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 1; act_sel_in[4] = 1; act_sel_in[5] = 4; act_sel_in[6] = 0; act_sel_in[7] = 3; act_sel_in[8] = 3; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 0; act_sel_in[12] = 1; act_sel_in[13] = 1; act_sel_in[14] = 0; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=4; act_sel_in[0] = 4; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 3; act_sel_in[4] = 4; act_sel_in[5] = 4; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 3; act_sel_in[9] = 0; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 0; act_sel_in[13] = 4; act_sel_in[14] = 3; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=3; act_sel_in[0] = 4; act_sel_in[1] = 0; act_sel_in[2] = 1; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 4; act_sel_in[6] = 0; act_sel_in[7] = 4; act_sel_in[8] = 4; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 1; act_sel_in[12] = 0; act_sel_in[13] = 0; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=2; act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 2; act_sel_in[3] = 3; act_sel_in[4] = 0; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 4; act_sel_in[9] = 3; act_sel_in[10] = 3; act_sel_in[11] = 3; act_sel_in[12] = 4; act_sel_in[13] = 1; act_sel_in[14] = 3; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 1; act_sel_in[5] = 0; act_sel_in[6] = 1; act_sel_in[7] = 1; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 0; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 1; act_sel_in[1] = 1; act_sel_in[2] = 4; act_sel_in[3] = 4; act_sel_in[4] = 0; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 1; act_sel_in[9] = 1; act_sel_in[10] = 1; act_sel_in[11] = 3; act_sel_in[12] = 1; act_sel_in[13] = 3; act_sel_in[14] = 1; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 


    #1 is_msb=1; column_idx=7; act_in[0] = -32; act_in[1] = -72; act_in[2] = 15; act_in[3] = -61; act_in[4] = 1; act_in[5] = 37; act_in[6] = 92; act_in[7] = -123; act_in[8] = 5; act_in[9] = 113; act_in[10] = 69; act_in[11] = 97; act_in[12] = -26; act_in[13] = -62; act_in[14] = 62; act_in[15] = 114; act_in[16] = 96; act_in[17] = 6; act_in[18] = 124; act_in[19] = -101; act_in[20] = 92; act_in[21] = -99; act_in[22] = 60; act_in[23] = 125; act_in[24] = -51; act_in[25] = 121; act_in[26] = 75; act_in[27] = 118; act_in[28] = 60; act_in[29] = -74; act_in[30] = 98; act_in[31] = -37; 
    act_sel_in[0] = 3; act_sel_in[1] = 3; act_sel_in[2] = 4; act_sel_in[3] = 1; act_sel_in[4] = 0; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 1; act_sel_in[9] = 0; act_sel_in[10] = 2; act_sel_in[11] = 2; act_sel_in[12] = 0; act_sel_in[13] = 2; act_sel_in[14] = 1; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 1; act_sel_in[3] = 3; act_sel_in[4] = 0; act_sel_in[5] = 1; act_sel_in[6] = 2; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 1; act_sel_in[11] = 4; act_sel_in[12] = 4; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=5; act_sel_in[0] = 1; act_sel_in[1] = 1; act_sel_in[2] = 2; act_sel_in[3] = 3; act_sel_in[4] = 3; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 4; act_sel_in[13] = 3; act_sel_in[14] = 3; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=4; act_sel_in[0] = 1; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 0; act_sel_in[5] = 2; act_sel_in[6] = 3; act_sel_in[7] = 0; act_sel_in[8] = 3; act_sel_in[9] = 0; act_sel_in[10] = 2; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 2; act_sel_in[3] = 1; act_sel_in[4] = 3; act_sel_in[5] = 0; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 4; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 3; act_sel_in[14] = 4; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=2; act_sel_in[0] = 0; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 3; act_sel_in[8] = 1; act_sel_in[9] = 4; act_sel_in[10] = 3; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 4; act_sel_in[14] = 1; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=1; act_sel_in[0] = 2; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 2; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 2; act_sel_in[7] = 0; act_sel_in[8] = 3; act_sel_in[9] = 2; act_sel_in[10] = 1; act_sel_in[11] = 0; act_sel_in[12] = 3; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=0; act_sel_in[0] = 2; act_sel_in[1] = 0; act_sel_in[2] = 0; act_sel_in[3] = 2; act_sel_in[4] = 2; act_sel_in[5] = 1; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 1; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 


    #1 is_msb=1; column_idx=7; act_in[0] = 32; act_in[1] = 81; act_in[2] = -66; act_in[3] = 98; act_in[4] = 7; act_in[5] = 62; act_in[6] = -54; act_in[7] = -118; act_in[8] = -86; act_in[9] = -18; act_in[10] = -9; act_in[11] = 119; act_in[12] = 91; act_in[13] = 96; act_in[14] = -120; act_in[15] = 20; act_in[16] = -95; act_in[17] = -43; act_in[18] = -47; act_in[19] = 35; act_in[20] = 87; act_in[21] = -45; act_in[22] = -128; act_in[23] = 90; act_in[24] = -88; act_in[25] = -27; act_in[26] = -110; act_in[27] = 13; act_in[28] = 43; act_in[29] = -59; act_in[30] = 87; act_in[31] = -22; 
    act_sel_in[0] = 4; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 3; act_sel_in[4] = 3; act_sel_in[5] = 1; act_sel_in[6] = 2; act_sel_in[7] = 2; act_sel_in[8] = 3; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 0; act_sel_in[12] = 1; act_sel_in[13] = 2; act_sel_in[14] = 1; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 0; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 4; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 0; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=5; act_sel_in[0] = 1; act_sel_in[1] = 0; act_sel_in[2] = 2; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 1; act_sel_in[8] = 4; act_sel_in[9] = 2; act_sel_in[10] = 2; act_sel_in[11] = 3; act_sel_in[12] = 4; act_sel_in[13] = 3; act_sel_in[14] = 4; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=4; act_sel_in[0] = 4; act_sel_in[1] = 0; act_sel_in[2] = 4; act_sel_in[3] = 0; act_sel_in[4] = 0; act_sel_in[5] = 3; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 1; act_sel_in[9] = 2; act_sel_in[10] = 1; act_sel_in[11] = 3; act_sel_in[12] = 3; act_sel_in[13] = 3; act_sel_in[14] = 0; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=3; act_sel_in[0] = 1; act_sel_in[1] = 0; act_sel_in[2] = 2; act_sel_in[3] = 3; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 0; act_sel_in[9] = 2; act_sel_in[10] = 2; act_sel_in[11] = 1; act_sel_in[12] = 2; act_sel_in[13] = 1; act_sel_in[14] = 1; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=2; act_sel_in[0] = 1; act_sel_in[1] = 1; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 1; act_sel_in[5] = 0; act_sel_in[6] = 1; act_sel_in[7] = 1; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 3; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=1; act_sel_in[0] = 0; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 3; act_sel_in[12] = 2; act_sel_in[13] = 1; act_sel_in[14] = 3; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=0; act_sel_in[0] = 4; act_sel_in[1] = 0; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 0; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 1; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 4; act_sel_in[12] = 3; act_sel_in[13] = 0; act_sel_in[14] = 3; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 


    #1 is_msb=1; column_idx=7; act_in[0] = 78; act_in[1] = 76; act_in[2] = 5; act_in[3] = -62; act_in[4] = -1; act_in[5] = -54; act_in[6] = -59; act_in[7] = -63; act_in[8] = 118; act_in[9] = 85; act_in[10] = 42; act_in[11] = -105; act_in[12] = 115; act_in[13] = -77; act_in[14] = 84; act_in[15] = 4; act_in[16] = 76; act_in[17] = -100; act_in[18] = 108; act_in[19] = 69; act_in[20] = -40; act_in[21] = -68; act_in[22] = -32; act_in[23] = -89; act_in[24] = 9; act_in[25] = -47; act_in[26] = -100; act_in[27] = 28; act_in[28] = 76; act_in[29] = -81; act_in[30] = 102; act_in[31] = -85; 
    act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 1; act_sel_in[3] = 0; act_sel_in[4] = 2; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 4; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 3; act_sel_in[11] = 3; act_sel_in[12] = 2; act_sel_in[13] = 0; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 3; act_sel_in[4] = 2; act_sel_in[5] = 3; act_sel_in[6] = 2; act_sel_in[7] = 2; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 3; act_sel_in[11] = 0; act_sel_in[12] = 3; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=5; act_sel_in[0] = 0; act_sel_in[1] = 0; act_sel_in[2] = 1; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 0; act_sel_in[11] = 2; act_sel_in[12] = 4; act_sel_in[13] = 4; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=4; act_sel_in[0] = 4; act_sel_in[1] = 0; act_sel_in[2] = 0; act_sel_in[3] = 3; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 3; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 0; act_sel_in[13] = 0; act_sel_in[14] = 3; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=3; act_sel_in[0] = 4; act_sel_in[1] = 3; act_sel_in[2] = 3; act_sel_in[3] = 4; act_sel_in[4] = 2; act_sel_in[5] = 1; act_sel_in[6] = 2; act_sel_in[7] = 2; act_sel_in[8] = 3; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 3; act_sel_in[12] = 1; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=2; act_sel_in[0] = 1; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 3; act_sel_in[4] = 0; act_sel_in[5] = 3; act_sel_in[6] = 2; act_sel_in[7] = 2; act_sel_in[8] = 3; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 4; act_sel_in[14] = 1; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=1; act_sel_in[0] = 3; act_sel_in[1] = 2; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 2; act_sel_in[5] = 4; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 3; act_sel_in[9] = 0; act_sel_in[10] = 3; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 3; act_sel_in[14] = 3; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 4; act_sel_in[6] = 1; act_sel_in[7] = 3; act_sel_in[8] = 1; act_sel_in[9] = 0; act_sel_in[10] = 2; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 


    #1 is_msb=1; column_idx=7; act_in[0] = 103; act_in[1] = 45; act_in[2] = 28; act_in[3] = -95; act_in[4] = -85; act_in[5] = 105; act_in[6] = -5; act_in[7] = 2; act_in[8] = 26; act_in[9] = 66; act_in[10] = 64; act_in[11] = 45; act_in[12] = -66; act_in[13] = -38; act_in[14] = -3; act_in[15] = 51; act_in[16] = 109; act_in[17] = 126; act_in[18] = -20; act_in[19] = 106; act_in[20] = -41; act_in[21] = 24; act_in[22] = 36; act_in[23] = -55; act_in[24] = -65; act_in[25] = -23; act_in[26] = 32; act_in[27] = 97; act_in[28] = -124; act_in[29] = -59; act_in[30] = 30; act_in[31] = 52; 
    act_sel_in[0] = 1; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 0; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 0; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 1; act_sel_in[1] = 0; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 4; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 3; act_sel_in[9] = 0; act_sel_in[10] = 0; act_sel_in[11] = 2; act_sel_in[12] = 4; act_sel_in[13] = 0; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=5; act_sel_in[0] = 1; act_sel_in[1] = 0; act_sel_in[2] = 0; act_sel_in[3] = 2; act_sel_in[4] = 3; act_sel_in[5] = 0; act_sel_in[6] = 1; act_sel_in[7] = 4; act_sel_in[8] = 2; act_sel_in[9] = 0; act_sel_in[10] = 1; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=4; act_sel_in[0] = 4; act_sel_in[1] = 3; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 1; act_sel_in[8] = 4; act_sel_in[9] = 3; act_sel_in[10] = 0; act_sel_in[11] = 4; act_sel_in[12] = 1; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 2; act_sel_in[3] = 3; act_sel_in[4] = 0; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 4; act_sel_in[9] = 3; act_sel_in[10] = 2; act_sel_in[11] = 1; act_sel_in[12] = 0; act_sel_in[13] = 2; act_sel_in[14] = 3; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=2; act_sel_in[0] = 4; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 0; act_sel_in[4] = 4; act_sel_in[5] = 2; act_sel_in[6] = 0; act_sel_in[7] = 0; act_sel_in[8] = 2; act_sel_in[9] = 1; act_sel_in[10] = 3; act_sel_in[11] = 2; act_sel_in[12] = 4; act_sel_in[13] = 0; act_sel_in[14] = 0; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=1; act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 4; act_sel_in[6] = 3; act_sel_in[7] = 2; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 2; act_sel_in[11] = 1; act_sel_in[12] = 2; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 2; act_sel_in[3] = 1; act_sel_in[4] = 0; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 1; act_sel_in[9] = 0; act_sel_in[10] = 0; act_sel_in[11] = 4; act_sel_in[12] = 3; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 


    #1 is_msb=1; column_idx=7; act_in[0] = -3; act_in[1] = 97; act_in[2] = -51; act_in[3] = 14; act_in[4] = 35; act_in[5] = -12; act_in[6] = 110; act_in[7] = 42; act_in[8] = 89; act_in[9] = 52; act_in[10] = -42; act_in[11] = 82; act_in[12] = -100; act_in[13] = 79; act_in[14] = -123; act_in[15] = -7; act_in[16] = 95; act_in[17] = 43; act_in[18] = -104; act_in[19] = -60; act_in[20] = 120; act_in[21] = -21; act_in[22] = -66; act_in[23] = 91; act_in[24] = 93; act_in[25] = 109; act_in[26] = -11; act_in[27] = -39; act_in[28] = 99; act_in[29] = -7; act_in[30] = 82; act_in[31] = -39; 
    act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 4; act_sel_in[3] = 4; act_sel_in[4] = 3; act_sel_in[5] = 3; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 1; act_sel_in[11] = 1; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 0; act_sel_in[4] = 2; act_sel_in[5] = 3; act_sel_in[6] = 3; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 3; act_sel_in[10] = 3; act_sel_in[11] = 2; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 1; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=5; act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 2; act_sel_in[3] = 3; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 0; act_sel_in[7] = 0; act_sel_in[8] = 2; act_sel_in[9] = 0; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 2; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=4; act_sel_in[0] = 2; act_sel_in[1] = 4; act_sel_in[2] = 1; act_sel_in[3] = 0; act_sel_in[4] = 0; act_sel_in[5] = 3; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 1; act_sel_in[9] = 4; act_sel_in[10] = 0; act_sel_in[11] = 2; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 4; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 3; act_sel_in[7] = 1; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 3; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=2; act_sel_in[0] = 3; act_sel_in[1] = 1; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 3; act_sel_in[5] = 0; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 3; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=1; act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 3; act_sel_in[3] = 4; act_sel_in[4] = 3; act_sel_in[5] = 0; act_sel_in[6] = 0; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 4; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 2; act_sel_in[1] = 0; act_sel_in[2] = 3; act_sel_in[3] = 2; act_sel_in[4] = 3; act_sel_in[5] = 4; act_sel_in[6] = 1; act_sel_in[7] = 4; act_sel_in[8] = 1; act_sel_in[9] = 3; act_sel_in[10] = 0; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 


    #1 is_msb=1; column_idx=7; act_in[0] = -98; act_in[1] = 63; act_in[2] = 44; act_in[3] = -117; act_in[4] = -25; act_in[5] = -98; act_in[6] = -91; act_in[7] = -38; act_in[8] = 120; act_in[9] = -78; act_in[10] = 21; act_in[11] = 125; act_in[12] = 15; act_in[13] = 112; act_in[14] = 119; act_in[15] = -18; act_in[16] = -70; act_in[17] = -112; act_in[18] = -101; act_in[19] = -23; act_in[20] = 120; act_in[21] = 101; act_in[22] = -89; act_in[23] = -48; act_in[24] = 53; act_in[25] = 26; act_in[26] = 123; act_in[27] = 5; act_in[28] = -66; act_in[29] = -43; act_in[30] = -33; act_in[31] = -83; 
    act_sel_in[0] = 1; act_sel_in[1] = 1; act_sel_in[2] = 2; act_sel_in[3] = 2; act_sel_in[4] = 0; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 4; act_sel_in[9] = 0; act_sel_in[10] = 1; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 2; act_sel_in[1] = 0; act_sel_in[2] = 0; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 4; act_sel_in[6] = 3; act_sel_in[7] = 1; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 0; act_sel_in[13] = 0; act_sel_in[14] = 0; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=5; act_sel_in[0] = 2; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 0; act_sel_in[5] = 1; act_sel_in[6] = 4; act_sel_in[7] = 1; act_sel_in[8] = 2; act_sel_in[9] = 1; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 1; act_sel_in[14] = 0; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=4; act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 3; act_sel_in[5] = 4; act_sel_in[6] = 4; act_sel_in[7] = 3; act_sel_in[8] = 2; act_sel_in[9] = 3; act_sel_in[10] = 4; act_sel_in[11] = 3; act_sel_in[12] = 3; act_sel_in[13] = 3; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 1; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 2; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 2; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=2; act_sel_in[0] = 2; act_sel_in[1] = 3; act_sel_in[2] = 0; act_sel_in[3] = 2; act_sel_in[4] = 3; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 2; act_sel_in[8] = 2; act_sel_in[9] = 2; act_sel_in[10] = 0; act_sel_in[11] = 4; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 2; act_sel_in[3] = 3; act_sel_in[4] = 4; act_sel_in[5] = 4; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 3; act_sel_in[9] = 2; act_sel_in[10] = 4; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 2; act_sel_in[14] = 3; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=0; act_sel_in[0] = 4; act_sel_in[1] = 4; act_sel_in[2] = 3; act_sel_in[3] = 0; act_sel_in[4] = 1; act_sel_in[5] = 1; act_sel_in[6] = 0; act_sel_in[7] = 3; act_sel_in[8] = 1; act_sel_in[9] = 4; act_sel_in[10] = 4; act_sel_in[11] = 1; act_sel_in[12] = 4; act_sel_in[13] = 0; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 


    #1 is_msb=1; column_idx=7; act_in[0] = 92; act_in[1] = 69; act_in[2] = 97; act_in[3] = -32; act_in[4] = -8; act_in[5] = 11; act_in[6] = -64; act_in[7] = 77; act_in[8] = -40; act_in[9] = 100; act_in[10] = 46; act_in[11] = -20; act_in[12] = 38; act_in[13] = 111; act_in[14] = 23; act_in[15] = 80; act_in[16] = -117; act_in[17] = 56; act_in[18] = -53; act_in[19] = -103; act_in[20] = -95; act_in[21] = 113; act_in[22] = -127; act_in[23] = -48; act_in[24] = -31; act_in[25] = 58; act_in[26] = 65; act_in[27] = -70; act_in[28] = 123; act_in[29] = -20; act_in[30] = 9; act_in[31] = -72; 
    act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 1; act_sel_in[3] = 0; act_sel_in[4] = 0; act_sel_in[5] = 1; act_sel_in[6] = 0; act_sel_in[7] = 2; act_sel_in[8] = 0; act_sel_in[9] = 2; act_sel_in[10] = 1; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 2; act_sel_in[1] = 3; act_sel_in[2] = 0; act_sel_in[3] = 1; act_sel_in[4] = 4; act_sel_in[5] = 1; act_sel_in[6] = 1; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 4; act_sel_in[10] = 4; act_sel_in[11] = 2; act_sel_in[12] = 3; act_sel_in[13] = 3; act_sel_in[14] = 4; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=5; act_sel_in[0] = 3; act_sel_in[1] = 2; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 3; act_sel_in[9] = 2; act_sel_in[10] = 3; act_sel_in[11] = 4; act_sel_in[12] = 3; act_sel_in[13] = 0; act_sel_in[14] = 0; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=4; act_sel_in[0] = 4; act_sel_in[1] = 1; act_sel_in[2] = 2; act_sel_in[3] = 1; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=3; act_sel_in[0] = 1; act_sel_in[1] = 1; act_sel_in[2] = 2; act_sel_in[3] = 3; act_sel_in[4] = 1; act_sel_in[5] = 0; act_sel_in[6] = 2; act_sel_in[7] = 4; act_sel_in[8] = 0; act_sel_in[9] = 1; act_sel_in[10] = 3; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=2; act_sel_in[0] = 0; act_sel_in[1] = 4; act_sel_in[2] = 1; act_sel_in[3] = 0; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 0; act_sel_in[7] = 1; act_sel_in[8] = 0; act_sel_in[9] = 2; act_sel_in[10] = 3; act_sel_in[11] = 4; act_sel_in[12] = 3; act_sel_in[13] = 0; act_sel_in[14] = 1; act_sel_in[15] = 1; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 0; act_sel_in[1] = 0; act_sel_in[2] = 3; act_sel_in[3] = 4; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 2; act_sel_in[9] = 3; act_sel_in[10] = 4; act_sel_in[11] = 0; act_sel_in[12] = 0; act_sel_in[13] = 4; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 4; act_sel_in[1] = 1; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 1; act_sel_in[5] = 3; act_sel_in[6] = 0; act_sel_in[7] = 3; act_sel_in[8] = 3; act_sel_in[9] = 0; act_sel_in[10] = 3; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 3; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 


    #1 is_msb=1; column_idx=7; act_in[0] = -31; act_in[1] = -121; act_in[2] = 16; act_in[3] = -112; act_in[4] = 46; act_in[5] = -78; act_in[6] = -127; act_in[7] = 57; act_in[8] = -56; act_in[9] = 34; act_in[10] = 52; act_in[11] = -38; act_in[12] = -29; act_in[13] = 107; act_in[14] = 96; act_in[15] = -51; act_in[16] = 30; act_in[17] = 59; act_in[18] = 84; act_in[19] = -97; act_in[20] = -87; act_in[21] = 36; act_in[22] = 29; act_in[23] = 123; act_in[24] = -102; act_in[25] = 87; act_in[26] = 54; act_in[27] = -4; act_in[28] = -11; act_in[29] = 90; act_in[30] = -64; act_in[31] = -72; 
    act_sel_in[0] = 1; act_sel_in[1] = 4; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 0; act_sel_in[5] = 0; act_sel_in[6] = 4; act_sel_in[7] = 4; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 3; act_sel_in[14] = 1; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 4; act_sel_in[1] = 0; act_sel_in[2] = 2; act_sel_in[3] = 4; act_sel_in[4] = 1; act_sel_in[5] = 4; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 1; act_sel_in[9] = 3; act_sel_in[10] = 0; act_sel_in[11] = 4; act_sel_in[12] = 3; act_sel_in[13] = 1; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=5; act_sel_in[0] = 1; act_sel_in[1] = 4; act_sel_in[2] = 4; act_sel_in[3] = 1; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 3; act_sel_in[8] = 3; act_sel_in[9] = 2; act_sel_in[10] = 3; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 0; act_sel_in[14] = 3; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=4; act_sel_in[0] = 3; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 0; act_sel_in[4] = 4; act_sel_in[5] = 4; act_sel_in[6] = 0; act_sel_in[7] = 4; act_sel_in[8] = 4; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 0; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 0; act_sel_in[4] = 0; act_sel_in[5] = 3; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 3; act_sel_in[9] = 4; act_sel_in[10] = 4; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 4; act_sel_in[14] = 3; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=2; act_sel_in[0] = 2; act_sel_in[1] = 0; act_sel_in[2] = 1; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 0; act_sel_in[7] = 0; act_sel_in[8] = 1; act_sel_in[9] = 1; act_sel_in[10] = 2; act_sel_in[11] = 1; act_sel_in[12] = 3; act_sel_in[13] = 3; act_sel_in[14] = 1; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=1; act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 2; act_sel_in[5] = 2; act_sel_in[6] = 0; act_sel_in[7] = 0; act_sel_in[8] = 4; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 2; act_sel_in[12] = 1; act_sel_in[13] = 0; act_sel_in[14] = 3; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 0; act_sel_in[1] = 3; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 3; act_sel_in[6] = 0; act_sel_in[7] = 3; act_sel_in[8] = 1; act_sel_in[9] = 0; act_sel_in[10] = 2; act_sel_in[11] = 2; act_sel_in[12] = 2; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 


    #1 is_msb=1; column_idx=7; act_in[0] = 72; act_in[1] = 41; act_in[2] = -43; act_in[3] = -79; act_in[4] = 121; act_in[5] = 17; act_in[6] = 119; act_in[7] = 46; act_in[8] = 72; act_in[9] = -7; act_in[10] = -25; act_in[11] = -73; act_in[12] = -91; act_in[13] = 73; act_in[14] = -105; act_in[15] = 73; act_in[16] = 107; act_in[17] = -98; act_in[18] = 49; act_in[19] = -101; act_in[20] = 101; act_in[21] = -84; act_in[22] = -84; act_in[23] = 50; act_in[24] = 84; act_in[25] = -17; act_in[26] = -64; act_in[27] = 50; act_in[28] = 9; act_in[29] = -13; act_in[30] = 0; act_in[31] = -12; 
    act_sel_in[0] = 1; act_sel_in[1] = 1; act_sel_in[2] = 4; act_sel_in[3] = 2; act_sel_in[4] = 3; act_sel_in[5] = 4; act_sel_in[6] = 2; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 3; act_sel_in[10] = 3; act_sel_in[11] = 3; act_sel_in[12] = 4; act_sel_in[13] = 4; act_sel_in[14] = 2; act_sel_in[15] = 3; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 4; act_sel_in[1] = 1; act_sel_in[2] = 3; act_sel_in[3] = 2; act_sel_in[4] = 4; act_sel_in[5] = 4; act_sel_in[6] = 4; act_sel_in[7] = 4; act_sel_in[8] = 3; act_sel_in[9] = 3; act_sel_in[10] = 2; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 3; act_sel_in[14] = 0; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=5; act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 0; act_sel_in[7] = 1; act_sel_in[8] = 2; act_sel_in[9] = 4; act_sel_in[10] = 0; act_sel_in[11] = 3; act_sel_in[12] = 0; act_sel_in[13] = 1; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 column_idx=4; act_sel_in[0] = 1; act_sel_in[1] = 3; act_sel_in[2] = 3; act_sel_in[3] = 3; act_sel_in[4] = 3; act_sel_in[5] = 1; act_sel_in[6] = 3; act_sel_in[7] = 1; act_sel_in[8] = 4; act_sel_in[9] = 2; act_sel_in[10] = 1; act_sel_in[11] = 1; act_sel_in[12] = 2; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=3; act_sel_in[0] = 3; act_sel_in[1] = 1; act_sel_in[2] = 4; act_sel_in[3] = 3; act_sel_in[4] = 4; act_sel_in[5] = 4; act_sel_in[6] = 1; act_sel_in[7] = 3; act_sel_in[8] = 3; act_sel_in[9] = 2; act_sel_in[10] = 3; act_sel_in[11] = 3; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 3; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=2; act_sel_in[0] = 2; act_sel_in[1] = 3; act_sel_in[2] = 3; act_sel_in[3] = 1; act_sel_in[4] = 0; act_sel_in[5] = 4; act_sel_in[6] = 4; act_sel_in[7] = 0; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 1; act_sel_in[11] = 3; act_sel_in[12] = 2; act_sel_in[13] = 1; act_sel_in[14] = 1; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=1; act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 3; act_sel_in[5] = 4; act_sel_in[6] = 4; act_sel_in[7] = 4; act_sel_in[8] = 1; act_sel_in[9] = 1; act_sel_in[10] = 0; act_sel_in[11] = 1; act_sel_in[12] = 1; act_sel_in[13] = 3; act_sel_in[14] = 0; act_sel_in[15] = 0; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=0; act_sel_in[0] = 4; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 2; act_sel_in[4] = 0; act_sel_in[5] = 3; act_sel_in[6] = 1; act_sel_in[7] = 4; act_sel_in[8] = 1; act_sel_in[9] = 2; act_sel_in[10] = 0; act_sel_in[11] = 3; act_sel_in[12] = 0; act_sel_in[13] = 4; act_sel_in[14] = 3; act_sel_in[15] = 2; act_val_in[0] = 1; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 


    #1 is_msb=1; column_idx=7; act_in[0] = 66; act_in[1] = 29; act_in[2] = 38; act_in[3] = -25; act_in[4] = -100; act_in[5] = -100; act_in[6] = 24; act_in[7] = -116; act_in[8] = -78; act_in[9] = -45; act_in[10] = -71; act_in[11] = -71; act_in[12] = -39; act_in[13] = -121; act_in[14] = -76; act_in[15] = -121; act_in[16] = -118; act_in[17] = -55; act_in[18] = -115; act_in[19] = -43; act_in[20] = 54; act_in[21] = -53; act_in[22] = -69; act_in[23] = 107; act_in[24] = 98; act_in[25] = -74; act_in[26] = 25; act_in[27] = -50; act_in[28] = -106; act_in[29] = 125; act_in[30] = -119; act_in[31] = -117; 
    act_sel_in[0] = 2; act_sel_in[1] = 1; act_sel_in[2] = 0; act_sel_in[3] = 2; act_sel_in[4] = 0; act_sel_in[5] = 4; act_sel_in[6] = 3; act_sel_in[7] = 3; act_sel_in[8] = 2; act_sel_in[9] = 3; act_sel_in[10] = 0; act_sel_in[11] = 4; act_sel_in[12] = 2; act_sel_in[13] = 4; act_sel_in[14] = 2; act_sel_in[15] = 1; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 1; 
    #1 is_msb=0; column_idx=6; act_sel_in[0] = 3; act_sel_in[1] = 1; act_sel_in[2] = 0; act_sel_in[3] = 4; act_sel_in[4] = 4; act_sel_in[5] = 0; act_sel_in[6] = 3; act_sel_in[7] = 1; act_sel_in[8] = 0; act_sel_in[9] = 2; act_sel_in[10] = 1; act_sel_in[11] = 3; act_sel_in[12] = 1; act_sel_in[13] = 1; act_sel_in[14] = 4; act_sel_in[15] = 2; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 1; is_skip_zero[1] = 0; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=5; act_sel_in[0] = 3; act_sel_in[1] = 2; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 3; act_sel_in[5] = 2; act_sel_in[6] = 4; act_sel_in[7] = 2; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 4; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 0; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 0; 
    #1 column_idx=4; act_sel_in[0] = 0; act_sel_in[1] = 2; act_sel_in[2] = 1; act_sel_in[3] = 1; act_sel_in[4] = 2; act_sel_in[5] = 3; act_sel_in[6] = 1; act_sel_in[7] = 1; act_sel_in[8] = 0; act_sel_in[9] = 0; act_sel_in[10] = 4; act_sel_in[11] = 3; act_sel_in[12] = 4; act_sel_in[13] = 4; act_sel_in[14] = 0; act_sel_in[15] = 3; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 0; act_val_in[4] = 1; act_val_in[5] = 1; act_val_in[6] = 1; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 1; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 0; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=3; act_sel_in[0] = 1; act_sel_in[1] = 2; act_sel_in[2] = 0; act_sel_in[3] = 0; act_sel_in[4] = 3; act_sel_in[5] = 0; act_sel_in[6] = 4; act_sel_in[7] = 0; act_sel_in[8] = 3; act_sel_in[9] = 2; act_sel_in[10] = 1; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 3; act_sel_in[14] = 3; act_sel_in[15] = 0; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 1; act_val_in[13] = 0; act_val_in[14] = 1; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=2; act_sel_in[0] = 0; act_sel_in[1] = 1; act_sel_in[2] = 3; act_sel_in[3] = 2; act_sel_in[4] = 0; act_sel_in[5] = 4; act_sel_in[6] = 1; act_sel_in[7] = 2; act_sel_in[8] = 0; act_sel_in[9] = 4; act_sel_in[10] = 2; act_sel_in[11] = 0; act_sel_in[12] = 2; act_sel_in[13] = 0; act_sel_in[14] = 4; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 0; act_val_in[2] = 0; act_val_in[3] = 1; act_val_in[4] = 1; act_val_in[5] = 0; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 0; is_skip_zero[0] = 0; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 
    #1 column_idx=1; act_sel_in[0] = 1; act_sel_in[1] = 1; act_sel_in[2] = 0; act_sel_in[3] = 3; act_sel_in[4] = 0; act_sel_in[5] = 2; act_sel_in[6] = 2; act_sel_in[7] = 4; act_sel_in[8] = 1; act_sel_in[9] = 2; act_sel_in[10] = 3; act_sel_in[11] = 4; act_sel_in[12] = 0; act_sel_in[13] = 2; act_sel_in[14] = 4; act_sel_in[15] = 4; act_val_in[0] = 0; act_val_in[1] = 1; act_val_in[2] = 0; act_val_in[3] = 0; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 1; act_val_in[8] = 0; act_val_in[9] = 0; act_val_in[10] = 1; act_val_in[11] = 0; act_val_in[12] = 0; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 0; is_skip_zero[3] = 0; 
    #1 column_idx=0; act_sel_in[0] = 1; act_sel_in[1] = 0; act_sel_in[2] = 1; act_sel_in[3] = 2; act_sel_in[4] = 1; act_sel_in[5] = 2; act_sel_in[6] = 1; act_sel_in[7] = 3; act_sel_in[8] = 0; act_sel_in[9] = 4; act_sel_in[10] = 1; act_sel_in[11] = 0; act_sel_in[12] = 4; act_sel_in[13] = 2; act_sel_in[14] = 2; act_sel_in[15] = 4; act_val_in[0] = 1; act_val_in[1] = 1; act_val_in[2] = 1; act_val_in[3] = 1; act_val_in[4] = 0; act_val_in[5] = 1; act_val_in[6] = 0; act_val_in[7] = 0; act_val_in[8] = 1; act_val_in[9] = 1; act_val_in[10] = 0; act_val_in[11] = 1; act_val_in[12] = 1; act_val_in[13] = 1; act_val_in[14] = 0; act_val_in[15] = 1; is_skip_zero[0] = 1; is_skip_zero[1] = 1; is_skip_zero[2] = 1; is_skip_zero[3] = 1; 



    #15 $stop;
  end

  always #1 clk = ~clk;

endmodule

`endif